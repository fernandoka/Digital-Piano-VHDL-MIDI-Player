----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Fernando Candelario Herrero
-- 
-- Create Date: 14.12.2019 20:22:30
-- Design Name: 
-- Module Name: MyDummyDDR2 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.4
-- Additional Comments:
--					 		
--
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MyDummyDDR2 is
  Port ( 
        rst_n           :   in  std_logic;
        clk             :   in  std_logic;
		addr			:	in	std_logic_vector(22 downto 0);
		cen             :	in	std_logic; -- low to request a read
        rd              :	in	std_logic; -- One cycle low to request a read
        wr              :	in	std_logic; -- One cycle low to request a read
		ack			    :	out	std_logic; -- One cycle high to notify the reception of a new byte
		data_in         :   in std_logic_vector(15 downto 0);
		data_out		:	out	std_logic_vector(127 downto 0)
  );
-- Attributes for debug
--attribute   dont_touch    :   string;
--attribute   dont_touch  of  MidiRom  :   entity  is  "true";
end MyDummyDDR2;

architecture Behavioral of MyDummyDDR2 is
	constant	MAX_ROWS	:	natural	:= 18256;
	
	type romType	is array (0 to MAX_ROWS) of std_logic_vector (127 downto 0);

    -- bach_tocatta_fugue_d_minor.mid
	constant romRd : romType :=(
    0=>X"544d000102000100060000006468544d", 1=>X"ff00081802040458ff009c0000006b72", 2=>X"ff0259ff0060e3160351ff0001ff0259", 3=>X"a160e3160351ff0040420f0351ff0001", 4=>X"40c3c027090351ff011516050351ff7f", 
    5=>X"479860e3160351ff60b6b0710b0351ff", 6=>X"00a8c027090351ff19811516050351ff", 7=>X"88862a2c0a0351ff0098804f120351ff", 8=>X"81d8b8050351ff61ae36140d0351ff00", 9=>X"009c36140d0351ff0036140d0351ff1f", 
    10=>X"ff0140420f0351ff00a020a1070351ff", 11=>X"b1000079b1001d7400006b72544d002f", 12=>X"c1006407b100330ab100305bb1000040", 13=>X"0ab100305bb1000040b1000079b10000", 14=>X"91006f6e6169500503ff006407b10033", 
    15=>X"91000051910000459110424591004651", 16=>X"9100004f91000043911045439100464f", 17=>X"51ff00404b4c0351ff20524591004f51", 18=>X"0351ff000051910000459140404b4c03", 19=>X"9100444f912060e3160351ff0060e316", 
    20=>X"9100444d9100004f9100004391104243", 21=>X"91004a4c9100004d9100004191104a41", 22=>X"9100444a9100004c9100004091104940", 23=>X"910047499100004a9100003e9110473e", 24=>X"9100504a910000499100003d91204d3d", 
    25=>X"4c0351ff0081004a9100003e91404c3e", 26=>X"3991004445910060e3160351ff40404b", 27=>X"3791004c439100004591000039911046", 28=>X"39910051459100004391000037911047", 29=>X"40404b4c0351ff00404b4c0351ff204d", 
    30=>X"ff0060e3160351ff0000459100003991", 31=>X"3491203e3491004440912060e3160351", 32=>X"35912049359100504191000040910000", 33=>X"31912048319100463d91000041910000", 34=>X"3291404f3291004c3e9100003d910000", 
    35=>X"51ff00404b4c0351ff0081003e910000", 36=>X"160351ff0060e3160351ff40404b4c03", 37=>X"9100002d9110472d91004639910060e3", 38=>X"9100002b9110482b91004d3791000039", 39=>X"4b4c0351ff204d2d9100523991000037", 
    40=>X"00399100002d9140404b4c0351ff0040", 41=>X"912060e3160351ff0060e3160351ff00", 42=>X"910000379100002b9110442b91004537", 43=>X"91000035910000299110472991004835", 44=>X"91000034910000289110472891004834", 
    45=>X"91000032910000269110482691004d32", 46=>X"91000031910000259120492591004c31", 47=>X"408100329100002691404f2691005332", 48=>X"31910082553191008244269100002691", 49=>X"00824e37910000349100824c34910000", 
    50=>X"4e3d9100003a910082433a9100003791", 51=>X"91110040916f8156409100003d910082", 52=>X"91004931910051409100513d9100513a", 53=>X"00003d91000040912381493791004934", 54=>X"0000319100003491000037915d003a91", 
    55=>X"40403291004c379100473e9100473991", 56=>X"8153369100003491404a349100003791", 57=>X"00399100003e91000032910000369100", 58=>X"3d91000031914041319100413d914083", 59=>X"3e91000032912a453291004e3e910000", 
    60=>X"4091000034912b4a3491004f40910000", 61=>X"3d91000031912b4a319100433d910000", 62=>X"3e91000032912a4d3291004c3e910000", 63=>X"4091000034912b4f3491005040910000", 64=>X"3d91000031912b48319100443d910000", 
    65=>X"3e91000032912a4a329100503e910000", 66=>X"4091000034912b4e3491004f40910000", 67=>X"3d91000031912b45319100463d910000", 68=>X"3e9100003291404f3291004c3e910000", 69=>X"409100003491404e3491005040910000", 
    70=>X"4191000035912a4b3591005141910000", 71=>X"4391000037912b4d3791005843910000", 72=>X"4091000034912b4a3491004740910000", 73=>X"4191000035912a4e3591004c41910000", 74=>X"4391000037912b513791005243910000", 
    75=>X"4091000034912b483491003e40910000", 76=>X"4191000035912a503591005041910000", 77=>X"4391000037912b513791004f43910000", 78=>X"4091000034912b4a3491004640910000", 79=>X"419100003591404b3591005341910000", 
    80=>X"43910000379140523791005443910000", 81=>X"4591000039912a513991005245910000", 82=>X"469100003a912b483a91004e46910000", 83=>X"4391000037912b4c3791004443910000", 84=>X"4591000039912a523991004d45910000", 
    85=>X"469100003a912b4d3a91005346910000", 86=>X"4391000037912b4b3791003e43910000", 87=>X"4591000039912a4f3991005045910000", 88=>X"469100003a912b4d3a91005046910000", 89=>X"4391000037912b493791004643910000", 
    90=>X"459100003991404f3991004c45910000", 91=>X"40404b4c0351ff00404b4c0351ff0000", 92=>X"914083c027090351ff00c027090351ff", 93=>X"910000499100003d9140443d91004749", 94=>X"9100004a9100003e912a503e91004b4a", 
    95=>X"9100004c91000040912b53409100554c", 96=>X"910000499100003d912b473d91004649", 97=>X"9100004a9100003e912a4c3e9100544a", 98=>X"9100004c91000040912b4e409100534c", 99=>X"910000499100003d912b4a3d91004449", 
    100=>X"9100004a9100003e912a4c3e9100504a", 101=>X"9100004c91000040912b51409100524c", 102=>X"910000499100003d912b463d91004349", 103=>X"9100004a9100003e91404f3e9100504a", 104=>X"9100004c91000040914050409100564c", 
    105=>X"9100004d91000041912a52419100524d", 106=>X"9100004f91000043912b504391004f4f", 107=>X"9100004c91000040912b4b409100484c", 108=>X"9100004d91000041912a514191004d4d", 109=>X"9100004f91000043912b4f439100514f", 
    110=>X"9100004c91000040912b45409100444c", 111=>X"9100004d91000041912a4f419100504d", 112=>X"9100004f91000043912b514391004d4f", 113=>X"9100004c91000040912b4b409100454c", 114=>X"9100004d910000419140514191004e4d", 
    115=>X"9100004f9100004391404a439100514f", 116=>X"9100005191000045912a514591005251", 117=>X"9100005291000046912b4c4691005152", 118=>X"9100004f91000043912b47439100434f", 119=>X"9100005191000045912a4d4591005251", 
    120=>X"9100005291000046912b524691004d52", 121=>X"9100004f91000043912b46439100484f", 122=>X"9100005191000045912a544591004a51", 123=>X"9100005291000046912b4c4691005052", 124=>X"9100004f91000043912b48439100464f", 
    125=>X"00840051910000459140514591004e51", 126=>X"00005191000045914040459100425191", 127=>X"00004f91000043912a49439100454f91", 128=>X"00005291000046912b524691004f5291", 129=>X"00004c91000040912b464091003c4c91", 
    130=>X"00004f91000043912a50439100524f91", 131=>X"00005291000046912b56469100525291", 132=>X"00004c91000040912b43409100464c91", 133=>X"00004d91000041912a504191004e4d91", 134=>X"00005191000045912b52459100525191", 
    135=>X"00004a9100003e912b453e91003f4a91", 136=>X"00004d91000041912a55419100514d91", 137=>X"00005191000045912b56459100555191", 138=>X"00004a9100003e912b3e3e91003f4a91", 139=>X"00004c91000040912a4b409100534c91", 
    140=>X"00004f91000043912b4f439100544f91", 141=>X"0000489100003c912b403c91003e4891", 142=>X"00004c91000040912a57409100524c91", 143=>X"00004f91000043912b56439100544f91", 144=>X"0000489100003c912b413c91003f4891", 
    145=>X"00004a9100003e912a4d3e91004d4a91", 146=>X"00004d91000041912b54419100514d91", 147=>X"0000469100003a912b483a9100414691", 148=>X"00004a9100003e912a563e91004d4a91", 149=>X"00004d91000041912b53419100534d91", 
    150=>X"0000469100003a912b463a9100414691", 151=>X"0000489100003c912a523c9100504891", 152=>X"00004c91000040912b59409100554c91", 153=>X"00004591000039912b453991003d4591", 154=>X"0000489100003c912a513c9100514891", 
    155=>X"00004c91000040912b55409100544c91", 156=>X"00004591000039912b4b399100424591", 157=>X"0000469100003a912a513a91004d4691", 158=>X"00004a9100003e912b533e9100514a91", 159=>X"00004391000037912b423791003e4391", 
    160=>X"0000469100003a912a493a9100504691", 161=>X"00004a9100003e912b513e9100544a91", 162=>X"00004391000037912b46379100414391", 163=>X"00004591000039912a4a399100504591", 164=>X"0000489100003c912b563c9100544891", 
    165=>X"00004191000035912b473591003b4191", 166=>X"00004591000039912a4f399100534591", 167=>X"0000489100003c912b543c9100554891", 168=>X"00004191000035912b47359100424191", 169=>X"00004391000037912a4d379100514391", 
    170=>X"0000469100003a912b483a9100504691", 171=>X"00004091000034912b43349100404091", 172=>X"00004391000037912a4e379100504391", 173=>X"0000469100003a912b513a9100504691", 174=>X"00004091000034912b473491003f4091", 
    175=>X"00004191000035912a4b3591004a4191", 176=>X"00004591000039912b53399100564591", 177=>X"00003e91000032912b423291003e3e91", 178=>X"00004191000035912a4c3591004f4191", 179=>X"00004591000039912b51399100554591", 
    180=>X"00003e91000032912b463291003d3e91", 181=>X"00004091000034912a4e3491004c4091", 182=>X"00004391000037912b513791004f4391", 183=>X"00003d91000031912b443191003f3d91", 184=>X"00004091000034912a51349100514091", 
    185=>X"00004391000037912b50379100554391", 186=>X"00003d91000031912b4b319100403d91", 187=>X"4243910042409100423d910082452691", 188=>X"58349100583191007f40b10042469100", 189=>X"379100003a910084583a910058379100", 
    190=>X"43910000269100003191000034910000", 191=>X"4691200040b100003d91000040910000", 192=>X"4391204a439100004591204745910000", 193=>X"40912043409100004191204541910000", 194=>X"3d9120453d9100003e9120463e910000", 
    195=>X"3d9140533d9100003b9120493b910000", 196=>X"3d9140533d9100003991404739910000", 197=>X"43912059439100004091205340910000", 198=>X"41911c474191060043911e4543910000", 199=>X"419118404191050043911a4543910500", 
    200=>X"4191164241910a0043911a4243910900", 201=>X"3e91004e419100004091404640910100", 202=>X"ff408142329100423991004235910044", 203=>X"00329140404b4c0351ff00404b4c0351", 204=>X"00419100003e91000035910000399100", 
    205=>X"4081b0710b0351ff00b0710b0351ff00", 206=>X"2044459120574a910000459140464591", 207=>X"204945910000459120534c9100004a91", 208=>X"204a45910000459120514d9100004c91", 209=>X"204b45910000459120444a9100004d91", 
    210=>X"2050459100004591204d4c9100004a91", 211=>X"204f459100004591204f4d9100004c91", 212=>X"204f45910000459120514f9100004d91", 213=>X"205245910000459120474c9100004f91", 214=>X"2043459120534d9100004c9100004591", 
    215=>X"204945910000459120524f9100004d91", 216=>X"204e4591000045912051519100004f91", 217=>X"204745910000459120424d9100005191", 218=>X"204b459100004591204e4f9100004d91", 219=>X"204d4591000045912057519100004f91", 
    220=>X"2046459100004591204f529100005191", 221=>X"204c45910000459120474f9100005291", 222=>X"204f459100004591204d519100004f91", 223=>X"204b45910000459120444d9100005191", 224=>X"204b459100004591204e4f9100004d91", 
    225=>X"204d45910000459120464c9100004f91", 226=>X"204d459100004591204d4d9100004c91", 227=>X"205145910000459120454a9100004d91", 228=>X"204a45910000459120524c9100004a91", 229=>X"204c459100004591204d499100004c91", 
    230=>X"20424591204f4a910000499100004591", 231=>X"204a4591000045912043459100004a91", 232=>X"204c459100004591204c469100004591", 233=>X"204b4591000045912045439100004691", 234=>X"2049459100004591204d459100004391", 
    235=>X"204b4591000045912046419100004591", 236=>X"204f4591000045912050439100004191", 237=>X"204b4591000045912046409100004391", 238=>X"204d459100004591204d419100004091", 239=>X"204d45910000459120463e9100004191", 
    240=>X"204c4591000045912052409100003e91", 241=>X"204845910000459120493d9100004091", 242=>X"204f459100004591204f419100003d91", 243=>X"204945910000459120453e9100004191", 244=>X"20494591000045912052409100003e91", 
    245=>X"204f45910000459120423d9100004091", 246=>X"2046459120523e9100003d9100004591", 247=>X"20484591000045912040399100003e91", 248=>X"2047459100004591204e3a9100003991", 249=>X"2048459100004591204a379100003a91", 
    250=>X"204b4591000045912049399100003791", 251=>X"20484591000045912048359100003991", 252=>X"204e459100004591204c379100003591", 253=>X"204f4591000045912051349100003791", 254=>X"2049459100004591204f359100003491", 
    255=>X"2048459100004591204c329100003591", 256=>X"204b4591000045912050379100003291", 257=>X"204d4591000045912046349100003791", 258=>X"204a459100004591204b359100003491", 259=>X"2049459100004591204b329100003591", 
    260=>X"204e459100004591204b349100003291", 261=>X"20514591000045912048319100003491", 262=>X"00329100814a32910000319100004591", 263=>X"0041912044419100003e9120453e9100", 264=>X"00419120434191000046912051469100", 
    265=>X"0040912044409100003c9120433c9100", 266=>X"00409120424091000045912055459100", 267=>X"003e9120423e9100003a9120413a9100", 268=>X"003e9120453e91000043912053439100", 269=>X"003d9120523d91000039912047399100", 
    270=>X"00459120554591000040912042409100", 271=>X"45419100003e914045329100413e9100", 272=>X"00419100004691000032914045469100", 273=>X"00309100003991405139910051309100", 274=>X"00409100004591404445910044409100", 
    275=>X"002e9100003a9140463a9100462e9100", 276=>X"003e91000043914045439100453e9100", 277=>X"452d9100453d91005045910050409100", 278=>X"3d9100002d9100003491008145349100", 279=>X"3e9120563e9100004091000045910000", 
    280=>X"4691205e469100004191204e41910000", 281=>X"3c9120493c9100004191204d41910000", 282=>X"45912060459100004091204a40910000", 283=>X"3a91204c3a9100004091204e40910000", 284=>X"43912061439100003e91204c3e910000", 
    285=>X"39912050399100003e91204c3e910000", 286=>X"4091204a409100003d91205c3d910000", 287=>X"3291004e3e9100004591205e45910000", 288=>X"3291404946910049419100003e91404b", 289=>X"39910052309100004191000046910000", 
    290=>X"45910046409100003091000039914052", 291=>X"3a91004b2e9100004091000045914046", 292=>X"439100493e9100002e9100003a91404b", 293=>X"45910055409100003e91000043914049", 294=>X"9100824a3491004a2d91004b3d910055", 
    295=>X"912000409100003d9100002d91000034", 296=>X"91204a419100004391204a4391000045", 297=>X"91204e3e9100004091204d4091000041", 298=>X"9120523b9100003d91204c3d9100003e", 299=>X"91204d399100003d9120593d9100003b", 
    300=>X"91205a3d9100003b9120553b91000039", 301=>X"91204b409100003e91205a3e9100003d", 302=>X"91205843910000419120584191000040", 303=>X"91204b43910000459120574591000043", 304=>X"91204e409100004191204d4191000043", 
    305=>X"91204a3e910000419120534191000040", 306=>X"91205a4591000041912058419100003e", 307=>X"91205c4a910000499120604991000045", 308=>X"9120564791000045912048459100004a", 309=>X"91205b4a910000499120564991000047", 
    310=>X"9110564d9100004c91205a4c9100004a", 311=>X"91205b519100004f9110564f9100004d", 312=>X"004b4a910000529100815a5291000051", 313=>X"404d5291004d4d9100004a91404c3291", 314=>X"004a459100004d910000529100003291", 
    315=>X"404c5191004c4c910000459140523091", 316=>X"004b469100004c910000519100003091", 317=>X"404d4f91004d4a910000469140522e91", 318=>X"005a499100004a9100004f9100002e91", 319=>X"81522d91004c4091005a5191005a4c91", 
    320=>X"004c91000051910000409100002d9100", 321=>X"4b4d9100004a9120644a910000499100", 322=>X"474d9100005291205f529100004d9120", 323=>X"574c91000048912045489100004d9120", 324=>X"494c91000051912061519100004c9120", 
    325=>X"484a9100004691204d469100004c9120", 326=>X"494a9100004f9120594f9100004a9120", 327=>X"60499100004591204e459100004a9120", 328=>X"5d519100004c91204a4c910000499120", 329=>X"004a91404a3291004f4a910000519120", 
    330=>X"00529100003291404d5291004d4d9100", 331=>X"00459140513091004a459100004d9100", 332=>X"00519100003091404c5191004c4c9100", 333=>X"00469140512e910048469100004c9100", 334=>X"004f9100002e91404c4f91004c4a9100", 
    335=>X"58519100584c910058499100004a9100", 336=>X"409100002d9100814f2d91004b409100", 337=>X"47910000499100004c91000051910000", 338=>X"2c910053419100533e9100533b910043", 339=>X"9100003e910000419100002c91008151", 
    340=>X"9100504091005249910000479100003b", 341=>X"404f47910000499140817e3991007e2b", 342=>X"000040910000479100002b9100003991", 343=>X"000049914060499100004591405d4591", 344=>X"00004f91205a4f9100004c91204a4c91", 
    345=>X"ff00005291405b529100404b4c0351ff", 346=>X"4f9100005191205651910060e3160351", 347=>X"4c9100004d9120514d9100004f91204f", 348=>X"4c9100004d9120534d9100004c912050", 349=>X"499100004a9120524a9100004c912050", 
    350=>X"489100004a91205a4a9100004991204b", 351=>X"4591000046912050469100004891204e", 352=>X"419100004391204d439100004591204f", 353=>X"3e910000409120544091000041912051", 354=>X"4691004e4c91004e499100003e912050", 
    355=>X"3d910063379100654391006540910061", 356=>X"91000043910000379100003d91008463", 357=>X"9100004991000040912a004c91000046", 358=>X"9100004c91000043912b7c439100594c", 359=>X"9100004991000040912b694091004b49", 
    360=>X"910000469100003d912a633d91004846", 361=>X"9100004991000040912b774091005849", 362=>X"910000469100003d912b683d91005046", 363=>X"9100004991000040912a794091005a49", 364=>X"9100004c91000043912b7c439100574c", 
    365=>X"9100004991000040912b634091004849", 366=>X"910000469100003d912a643d91004f46", 367=>X"9100004991000040912b754091005649", 368=>X"910000469100003d912b6d3d91004f46", 369=>X"9100004991000040912a784091005a49", 
    370=>X"9100004c91000043912b764391005e4c", 371=>X"9100004991000040912b674091004a49", 372=>X"910000469100003d912a643d91004a46", 373=>X"9100004991000040912b7e4091005749", 374=>X"910000469100003d912b653d91004d46", 
    375=>X"9100004991000040912a7a4091006049", 376=>X"9100004c91000043912b7b4391005c4c", 377=>X"9100004991000040912b6c4091004e49", 378=>X"910000469100003d912a673d91004c46", 379=>X"9100004991000040912b7c4091005e49", 
    380=>X"910000469100003d912b663d91004f46", 381=>X"910000439100003a912a6c3a91004c43", 382=>X"910000469100003d912b783d91005746", 383=>X"910000439100003a912b713a91004e43", 384=>X"9100004091000037912a673791004a40", 
    385=>X"910000439100003a912b753a91005a43", 386=>X"9100004091000037912b6b3791004d40", 387=>X"910000439100003a912a753a91005c43", 388=>X"910000469100003d912b7d3d91005646", 389=>X"910000439100003a912b6c3a91004d43", 
    390=>X"9100004091000037912a6b3791004640", 391=>X"910000439100003a912b763a91005c43", 392=>X"9100004091000037912b6b3791004b40", 393=>X"910000439100003a912a733a91005843", 394=>X"910000469100003d912b7d3d91005d46", 
    395=>X"910000439100003a912b6c3a91004d43", 396=>X"9100004091000037912a6b3791004c40", 397=>X"910000439100003a912b723a91005643", 398=>X"9100004091000037912b6e3791004c40", 399=>X"910000439100003a912a753a91005b43", 
    400=>X"910000469100003d912b7b3d91005b46", 401=>X"910000439100003a912b6f3a91005143", 402=>X"9100004091000037912a6e3791004940", 403=>X"910000439100003a912b763a91005843", 404=>X"9100004091000037912b6f3791004b40", 
    405=>X"9100003d91000034912a663491004c3d", 406=>X"9100004091000037912b743791005840", 407=>X"9100003d91000034912b6a3491004a3d", 408=>X"9100003a91000031912a6f319100513a", 409=>X"9100003d91000034912b773491005e3d", 
    410=>X"9100003a91000031912b6e319100543a", 411=>X"9100003d91000034912a753491005b3d", 412=>X"9100004091000037912b773791005b40", 413=>X"9100003d91000034912b6e3491004e3d", 414=>X"9100003a91000031912a6a3191004b3a", 
    415=>X"9100003d91000034912b76349100593d", 416=>X"9100003a91000031912b6c3191004c3a", 417=>X"9100003d91000034912a75349100583d", 418=>X"9100004091000037912b783791005a40", 419=>X"9100003d91000034912b693491004a3d", 
    420=>X"9100003a91000031912a68319100453a", 421=>X"9100003d91000034912b713491005b3d", 422=>X"9100003a91000031912b6c319100513a", 423=>X"9100003d91000034912a76349100593d", 424=>X"9100004091000037912b713791005c40", 
    425=>X"9100003d91000034912b733491004f3d", 426=>X"9100003a91000031912a70319100523a", 427=>X"9100003d91000034912b72349100593d", 428=>X"9100003a91000031912b6c3191004e3a", 429=>X"9100003d91000034912a703491005e3d", 
    430=>X"9100004091000037912b753791005b40", 431=>X"9100003d91000034912b703491004b3d", 432=>X"9100004091000037912a773791005740", 433=>X"910000439100003a912b703a91005c43", 434=>X"9100004091000037912b703791005340", 
    435=>X"9100003d91000034912a6b349100493d", 436=>X"9100004091000037912b723791005840", 437=>X"9100003d91000034912b723491004c3d", 438=>X"9100004091000037912a783791005e40", 439=>X"910000439100003a912b753a91005843", 
    440=>X"9100004091000037912b6c3791005040", 441=>X"9100003d91000034912a6e3491004c3d", 442=>X"9100004091000037912b773791005840", 443=>X"9100003d91000034912b693491004e3d", 444=>X"9100004091000037912a783791005840", 
    445=>X"910000439100003a912b763a91005f43", 446=>X"9100004091000037912b693791004b40", 447=>X"9100003d91000034912a6a3491004b3d", 448=>X"9100004091000037912b763791005740", 449=>X"9100003d91000034912b6d3491004e3d", 
    450=>X"9100004091000037912a773791005840", 451=>X"910000439100003a912b773a91005943", 452=>X"9100004091000037912b6e3791004940", 453=>X"9100004391000034912a6a3491005843", 454=>X"9100004691000037912b763791005646", 
    455=>X"9100004391000034912b6b3491004d43", 456=>X"9100004691000034912a723491005946", 457=>X"9100004391000037912b773791005243", 458=>X"9100004691000034912b6d3491005746", 459=>X"910000439100003a912a7e3a91004a43", 
    460=>X"910000469100003d912b7e3d91005b46", 461=>X"910000439100003a912b723a91005043", 462=>X"910000469100003a912a713a91005b46", 463=>X"910000439100003d912b7a3d91004a43", 464=>X"910000469100003a912b6f3a91005c46", 
    465=>X"9100004991000040912a7e4091005b49", 466=>X"910000469100003d912b6a3d91005246", 467=>X"9100004991000040912b7a4091005d49", 468=>X"9100004c9100003d912a6c3d91005c4c", 469=>X"9100004991000040912b744091005349", 
    470=>X"9100004c9100003d912b6a3d91005f4c", 471=>X"9100004991000040912a7b4091004a49", 472=>X"9100004c9100003d912b6a3d91005d4c", 473=>X"9100004991000040912b774091004a49", 474=>X"9100004c9100003d912a693d91005c4c", 
    475=>X"9100004991000040912b7a4091004c49", 476=>X"9100004c9100003d912b6c3d9100594c", 477=>X"910062519100624c9100624991006245", 478=>X"008265399100653791004a4091004a3d", 479=>X"00003d91000040910000379100003991", 
    480=>X"000045910000499100004c9100005191", 481=>X"0054519100544d9100544a9100544591", 482=>X"826a3991006a35910059419100593e91", 483=>X"003e9100004191000035910000399100", 484=>X"00459100004a9100004d910000519100", 
    485=>X"593e91004a4f91004a4a91004a469100", 486=>X"3e91000043910082713a910059439100", 487=>X"91008100469100004a9100004f910000", 488=>X"91406e379100003991406c399100003a", 489=>X"91004e4c91004e4991004e4591000037", 
    490=>X"4081773991004b4091004b3d91004e4f", 491=>X"00004091000034914069349100003991", 492=>X"0000499100004c9100004f9100003d91", 493=>X"406d3291000035914075359100004591", 494=>X"406f3191000034914077349100003291", 
    495=>X"40712f91000032914072329100003191", 496=>X"406a2d91000031914078319100002f91", 497=>X"406e2c9100002e9140772e9100002d91", 498=>X"004c459100002d9140772d9100002c91", 499=>X"00003991407e3991004e4091004c4991", 
    500=>X"005d4191000045910000499100004091", 501=>X"0072359100513e91005d4a91005d4591", 502=>X"003e9100003591000039910081723991", 503=>X"3e4191000041910000459100004a9100", 504=>X"329100816b3991006b329100563e9100", 
    505=>X"9100816f2d91004e4091000041910000", 506=>X"9100002d910000399140503d9100003e", 507=>X"9100503e910000409100003d91407037", 508=>X"00003791008168329100682691006639", 509=>X"000034914070349100003591406f3591", 
    510=>X"00269100003291000035910082743591", 511=>X"004591405e459140003e910000399100", 512=>X"004591406a459100004391405f439100", 513=>X"00459140694591000041914056419100", 514=>X"004591406d4591000040914056409100", 
    515=>X"0045914071459100003e9140503e9100", 516=>X"004591406c459100003d9140503d9100", 517=>X"004591406d459100003e9140523e9100", 518=>X"00459140684591000040914058409100", 519=>X"004591406d459100004191405a419100", 
    520=>X"00459140794591000039914051399100", 521=>X"004591407a459100003b91405a3b9100", 522=>X"0045914071459100003d9140523d9100", 523=>X"0045914074459100003e9140533e9100", 524=>X"004591406f459100003d91404f3d9100", 
    525=>X"0045914073459100003e9140563e9100", 526=>X"00459140694591000040914056409100", 527=>X"004a9100004191405b4a914059419100", 528=>X"694a9100004891406542910056489100", 529=>X"6343910056469100004a910000429140", 
    530=>X"004a9100004391406b4a910000469140", 531=>X"704a9100004591404d3c910055459100", 532=>X"5a3a910051439100004a9100003c9140", 533=>X"004a9100003a91406e4a910000439140", 534=>X"704a9100004291405d39910050429100", 
    535=>X"623a910051439100004a910000399140", 536=>X"004a9100003a91406f4a910000439140", 537=>X"6b4a910000459140673c910053459100", 538=>X"6c3e91005c469100004a9100003c9140", 539=>X"004a9100003e9140684a910000469140", 
    540=>X"754a9100003e91405d369100483e9100", 541=>X"613791004e409100004a910000369140", 542=>X"004a9100003791407b4a910000409140", 543=>X"734a9100004291406239910054429100", 544=>X"623a91004f439100004a910000399140", 
    545=>X"004a9100003a9140704a910000439140", 546=>X"724a9100004291405d3991004e429100", 547=>X"633a910052439100004a910000399140", 548=>X"004a9100003a9140734a910000439140", 549=>X"6a4a9100004591405f36910057459100", 
    550=>X"623791005b469100004a910000369140", 551=>X"00469100004391407d43910000379140", 552=>X"7c4391000037914059379100684a9100", 553=>X"5b3e91005b469100004a910000439140", 554=>X"00469100004391406c439100003e9140", 
    555=>X"72439100003e9140543e9100674a9100", 556=>X"4a3c9100674b9100004a910000439140", 557=>X"004b9100003f9140673f9100003c9140", 558=>X"693f9100003c9140593c91004f439100", 559=>X"5b3c9100704b910000439100003f9140", 
    560=>X"004b9100003f91406a3f9100003c9140", 561=>X"6b3f9100003c9140543c91004d439100", 562=>X"5d3c91006848910000439100003f9140", 563=>X"004891000041914073419100003c9140", 564=>X"6a419100003c91405a3c91005b459100", 
    565=>X"563c9100684891000045910000419140", 566=>X"00489100004191406f419100003c9140", 567=>X"6c419100003c9140563c910057459100", 568=>X"593a91006c4a91000045910000419140", 569=>X"004a9100003e91406a3e9100003a9140", 
    570=>X"6a3e9100003a91405d3a91004e419100", 571=>X"5c3a9100724a910000419100003e9140", 572=>X"004a9100003e91406a3e9100003a9140", 573=>X"693e9100003a9140603a91004e419100", 574=>X"623a91006746910000419100003e9140", 
    575=>X"00469100004091406f409100003a9140", 576=>X"6f409100003a91405b3a91005b439100", 577=>X"5f3a91006d4691000043910000409140", 578=>X"004691000040914070409100003a9140", 579=>X"72409100003a91405a3a91005c439100", 
    580=>X"5d3991006d4991000043910000409140", 581=>X"00499100003d9140693d910000399140", 582=>X"6a3d9100003991406339910051409100", 583=>X"5c3991007249910000409100003d9140", 584=>X"00499100003d9140723d910000399140", 
    585=>X"6b3d9100003991405e3991004b409100", 586=>X"593591006e45910000409100003d9140", 587=>X"00459100003e9140753e910000359140", 588=>X"7a3e910000359140583591005a419100", 589=>X"5e3591006a45910000419100003e9140", 
    590=>X"00459100003e9140783e910000359140", 591=>X"723e9100003591405a3591005c419100", 592=>X"5b3491006443910000419100003e9140", 593=>X"00439100003a9140693a910000349140", 594=>X"673a910000349140563491004e3d9100", 
    595=>X"5c34910071439100003d9100003a9140", 596=>X"00439100003a91406b3a910000349140", 597=>X"673a91000034914059349100573d9100", 598=>X"563291006b419100003d9100003a9140", 599=>X"00419100003991406839910000329140", 
    600=>X"63399100003291405c3291005b3e9100", 601=>X"5c32910066419100003e910000399140", 602=>X"00419100003991406939910000329140", 603=>X"6539910000329140593291005a3e9100", 604=>X"583491004a409100003e910000399140", 
    605=>X"0037914064379100003491010040913f", 606=>X"00349101003a913f5e3491004a3a9100", 607=>X"61349100604091000037914066379100", 608=>X"0037914065379100003491010040913f", 609=>X"00349101003a913f5d3491004b3a9100", 
    610=>X"61359100563991000037914065379100", 611=>X"00519100003991000035914055519140", 612=>X"004f9140623491005c3991005d4f9100", 613=>X"00519100003991000034914065519100", 614=>X"004d91405b3291005f399100584d9100", 
    615=>X"00519100003991000032914069519100", 616=>X"004c91406837910061399100554c9100", 617=>X"0051910000399100003791406c519100", 618=>X"004a91405e3591005f399100534a9100", 619=>X"00519100003991000035914074519100", 
    620=>X"004991405a3491006139910051499100", 621=>X"00519100003991000034914072519100", 622=>X"004a91406635910061399100514a9100", 623=>X"00519100003991000035914072519100", 624=>X"004c91405c31910063399100584c9100", 
    625=>X"00519100003991000031914068519100", 626=>X"004d91405f329100603991005c4d9100", 627=>X"00519100003991000032914069519100", 628=>X"004591405d3191006339910044459100", 629=>X"00519100003991000031914076519100", 
    630=>X"00479140633291005d3991004b479100", 631=>X"00519100003991000032914075519100", 632=>X"00499140603491006339910052499100", 633=>X"0051910000399100003491406f519100", 634=>X"004a91405f35910065399100524a9100", 
    635=>X"00519100003991000035914072519100", 636=>X"004991405e3491005d39910050499100", 637=>X"00519100003991000034914076519100", 638=>X"004a91406635910061399100524a9100", 639=>X"0051910000399100003591406f519100", 
    640=>X"004c91405d31910064399100564c9100", 641=>X"0051910000399100003191406c519100", 642=>X"004d914061329100613991005b4d9100", 643=>X"004c9140534c91000051914069519100", 644=>X"0051910000399100003291406d519100", 
    645=>X"004a914065359100703e9100534a9100", 646=>X"004891404d489100005191406e519100", 647=>X"00519100003e91000035914075519100", 648=>X"0046914063379100663e91004a469100", 649=>X"004891404c4891000051914077519100", 
    650=>X"00519100003e91000037914072519100", 651=>X"004f91406d4f9100004a9140534a9100", 652=>X"004f91406f4f9100004691404a469100", 653=>X"004c9140583091005c3c91005d4c9100", 654=>X"004a9140504a9100004f91406a4f9100", 
    655=>X"004f9100003c9100003091406c4f9100", 656=>X"004891406b349100623c910051489100", 657=>X"004691404f469100004f9140714f9100", 658=>X"004f9100003c910000349140764f9100", 659=>X"00459140643591005d3c91004e459100", 
    660=>X"0046914050469100004f9140764f9100", 661=>X"004f9100003c910000359140704f9100", 662=>X"004d91406d4d91000048914052489100", 663=>X"004d9140704d91000045914051459100", 664=>X"004a91405a2e9100573a91005a4a9100", 
    665=>X"0048914052489100004d9140694d9100", 666=>X"004d9100003a9100002e91406b4d9100", 667=>X"00469140653291005c3a910054469100", 668=>X"0045914051459100004d9140744d9100", 669=>X"004d9100003a9100003291406f4d9100", 
    670=>X"0043914065349100643a910052439100", 671=>X"0045914053459100004d9140764d9100", 672=>X"004d9100003a910000349140734d9100", 673=>X"004c9140724c91000046914055469100", 674=>X"004c91406f4c9100004391404f439100", 
    675=>X"00499140542d91005539910060499100", 676=>X"0046914054469100004c91406c4c9100", 677=>X"004c910000399100002d91406e4c9100", 678=>X"00459140653191006439910054459100", 679=>X"004391404e439100004c9140774c9100", 
    680=>X"004c91000039910000319140754c9100", 681=>X"0041914063329100623991004a419100", 682=>X"0043914052439100004c9140744c9100", 683=>X"004c91000039910000329140714c9100", 684=>X"004a91406e4a91000045914057459100", 
    685=>X"004191405a3591004b3e91004b419100", 686=>X"003e9100004a9100003591406f4a9100", 687=>X"00409140653a9100483d91004f409100", 688=>X"003d9100004c9100003a91407b4c9100", 689=>X"00409140623a9100513d910047409100", 
    690=>X"003d9100004c9100003a9140774c9100", 691=>X"0041914060399100593e91004e419100", 692=>X"003e9100004a910000399140744a9100", 693=>X"0041914065399100513e91004c419100", 694=>X"003e9100004a910000399140724a9100", 
    695=>X"00469140603791005e4091005c469100", 696=>X"004691405a469100004991406c499100", 697=>X"00409100004991000037914069499100", 698=>X"004a9140684a91000045914055459100", 699=>X"004191405a3991004f3e910050419100", 
    700=>X"003e9100004a910000399140734a9100", 701=>X"00409140633a91004c3d91004b409100", 702=>X"003d9100004c9100003a91407c4c9100", 703=>X"00409140663a91004e3d91004a409100", 704=>X"003d9100004c9100003a91407b4c9100", 
    705=>X"0041914060399100573e91004b419100", 706=>X"003e9100004a910000399140724a9100", 707=>X"0041914060399100593e91004e419100", 708=>X"003e9100004a9100003991406f4a9100", 709=>X"004a9140544a91405f38910057409100", 
    710=>X"00389140634a9100004991405b499100", 711=>X"004791405747910000409100004a9100", 712=>X"004991405d499100004a9140674a9100", 713=>X"4b45914064499100004791405a479100", 714=>X"51459100004391404d43910000459140", 
    715=>X"004091404c4091000049910000459140", 716=>X"004191404b419100004391405c439100", 717=>X"584a91405d419100004091404c409100", 718=>X"664a9100004991405a499100004a9140", 719=>X"4f3e91006b4d910000419100004a9140", 
    720=>X"60499100004a91405b4a9100004d9140", 721=>X"003e9100004791405a47910000499140", 722=>X"69459100003991404f39910066499100", 723=>X"5f459100004391405443910000459140", 724=>X"483d9100674c91000049910000459140", 
    725=>X"4f419100004391405c439100003d9140", 726=>X"59419100004091405440910000419140", 727=>X"5b4a9100004c9100003e9140573e9140", 728=>X"003e9140603e9100003d91405c3d9100", 729=>X"00399140583991005240910000419100", 
    730=>X"5a499100004a9100003991405f399100", 731=>X"0039914063399100003791405c379100", 732=>X"493e91005b4891000040910000499100", 733=>X"003e9140743e91000036914058369100", 734=>X"003d9140623d910064459100003e9100", 
    735=>X"5e46910000489100003e9140663e9100", 736=>X"00419140764191000037914057379100", 737=>X"003f9140603f91004e43910000459100", 738=>X"5d45910000469100003e91405a3e9100", 739=>X"0040914067409100003d91405a3d9100", 
    740=>X"003d91406d3d91000039914057399100", 741=>X"4c429100654591000045910000439100", 742=>X"003f91407e3f91000032914054329100", 743=>X"003c91405b3c9100003e9140653e9100", 744=>X"53419100584391000045910000429100", 
    745=>X"003e91406a3e9100003b9140603b9100", 746=>X"003b9140643b9100003791405d379100", 747=>X"4e3f9100604391000043910000419100", 748=>X"003e91407b3e91000030914057309100", 749=>X"003a9140603a9100003c91405f3c9100", 
    750=>X"003991405e3991005e42910000439100", 751=>X"00429100003f9100003c91406a3c9100", 752=>X"003691405c3691004e3e910068459100", 753=>X"60429100003e91000039914064399100", 754=>X"003c91407c3c91000032914053329100", 
    755=>X"62489100714b91000045910000429100", 756=>X"003991405d399100003a9140603a9100", 757=>X"003a9140623a91005d4a9100004b9100", 758=>X"4a46910000489100004591407c459100", 759=>X"4e45910000469100004391405b439100", 
    760=>X"004a910000459100004291405c429100", 761=>X"583a9100004391406243910051469100", 762=>X"504691005a4f910000469100003a9140", 763=>X"003791405c379100003991405c399100", 764=>X"00329140593291404c45910000469100", 
    765=>X"003091405c3091005a4e9100004f9100", 766=>X"00459100004e91000032914065329100", 767=>X"002e9140632e91005d4a9100634f9100", 768=>X"50489100004a91000032914062329100", 769=>X"0032914067329100002d91405d2d9100", 
    770=>X"5146910049469100004f910000489100", 771=>X"0032914066329100002b91405b2b9100", 772=>X"4e459100694a91000046910000469100", 773=>X"0032914067329100002a9140582a9100", 774=>X"544691005f4a9100004a910000459100", 
    775=>X"003291406c329100002b91405c2b9100", 776=>X"4b429100614a9100004a910000469100", 777=>X"0032914062329100002d9140632d9100", 778=>X"55439100644a9100004a910000429100", 779=>X"0032914065329100002e91405e2e9100", 
    780=>X"554291005f4a9100004a910000439100", 781=>X"003291406d3291000026914055269100", 782=>X"504391005e4a9100004a910000429100", 783=>X"00329140663291000028914059289100", 784=>X"56459100604a9100004a910000439100", 
    785=>X"0032914068329100002a91405c2a9100", 786=>X"574691005f4a9100004a910000459100", 787=>X"003291406e329100002b9140582b9100", 788=>X"51459100624a9100004a910000469100", 789=>X"003291406b329100002a9140552a9100", 
    790=>X"53469100604a9100004a910000459100", 791=>X"0032914069329100002b9140572b9100", 792=>X"4d429100604a9100004a910000469100", 793=>X"0032914067329100002d91405c2d9100", 794=>X"554391005f4a9100004a910000429100", 
    795=>X"004a9100004391406c3a91006c2e9100", 796=>X"004f910000469140594691006e4f9100", 797=>X"004d910000459140524591005e4d9100", 798=>X"002e9100003a914056469100684f9100", 799=>X"4e439100594c9100004f910000469100", 
    800=>X"59459100674d9100004c910000439140", 801=>X"4c4191005a4a9100004d910000459140", 802=>X"674c9100004a910000419140592f9100", 803=>X"004c910000439100002f914053439100", 804=>X"004091405e3091004d40910055489100", 
    805=>X"004891405f4891007451910000489100", 806=>X"0046914053469100594f910000519100", 807=>X"003091405e4891006b519100004f9100", 808=>X"4d459100544d91000051910000489100", 809=>X"5a469100644f9100004d910000459140", 
    810=>X"4d439100574c9100004f910000469140", 811=>X"664d9100004c91000043914056319100", 812=>X"004d910000459100003191405a459100", 813=>X"00419140643291004e419100574a9100", 814=>X"004a9140634a910075529100004a9100", 
    815=>X"00489140514891006151910000529100", 816=>X"00329140584a91006552910000519100", 817=>X"48469100584f910000529100004a9100", 818=>X"5548910064519100004f910000469140", 819=>X"47459100564d91000051910000489140", 
    820=>X"604f9100004d91000045914053329100", 821=>X"004f910000469100003291405b469100", 822=>X"004391405e3491004d4391005a4c9100", 823=>X"004c91405f4c910077549100004c9100", 824=>X"004a9140514a91006052910000549100", 
    825=>X"003491405d4c91006b54910000529100", 826=>X"494891005a51910000549100004c9100", 827=>X"594a9100635291000051910000489140", 828=>X"494691005a4f910000529100004a9140", 829=>X"69519100004f91000046914055349100", 
    830=>X"0051910000489100003491405a489100", 831=>X"004d9140623591004b459100574d9100", 832=>X"00459100004b9100003591405a4b9100", 833=>X"004a91405c2d91004c4191005e4a9100", 834=>X"0041910000489100002d914059489100", 
    835=>X"004691405d2e91005e4691006b4a9100", 836=>X"002e9140514591005d489100004a9100", 837=>X"50439100574691000048910000459100", 838=>X"5f459100004691000043914066329100", 839=>X"00459100004191000032914046419100", 
    840=>X"00439140582b91005743910064469100", 841=>X"004691405d4691006f4a910000469100", 842=>X"004391404b4391005d469100004a9100", 843=>X"002b91404c4191005a45910000469100", 844=>X"4f4091005c4391000045910000419100", 
    845=>X"58439100684691000043910000409140", 846=>X"4c4091005a4391000046910000439140", 847=>X"594191000043910000409140572e9100", 848=>X"5d40910000419100003e91404f3e9100", 849=>X"6641910000409100003c91404c3c9100", 
    850=>X"00419100003e9100002e9140583e9100", 851=>X"00409140612d91005e4091006a439100", 852=>X"002d91405d4191006a45910000439100", 853=>X"5b4391006a4691000045910000419100", 854=>X"002b91406d4a910000469140602b9100", 
    855=>X"4e4091005f48910000439100004a9100", 856=>X"003091405c4691000048914066309100", 857=>X"5b4191005d4591000040910000469100", 858=>X"003c91407d3c9100002991405e299100", 859=>X"003c9140653c9100003a9140623a9100", 
    860=>X"5d399100694891000045910000419100", 861=>X"00489100003c9140643c910000399140", 862=>X"673c910000379140613791005a469100", 863=>X"583591005d45910000469100003c9140", 864=>X"00459100003c91406d3c910000359140", 
    865=>X"743c9100003491405834910058439100", 866=>X"5d3591006545910000439100003c9140", 867=>X"00459100003c9140713c910000359140", 868=>X"6b3c9100003791406237910067469100", 869=>X"5c3991006848910000469100003c9140", 
    870=>X"00489100003c91406e3c910000399140", 871=>X"793c9100003091405630910050409100", 872=>X"583291006341910000409100003c9140", 873=>X"00419100003c9140763c910000329140", 874=>X"773c9100003491405934910069439100", 
    875=>X"5f3591006b45910000439100003c9140", 876=>X"00459100003c9140703c910000359140", 877=>X"763c9100003491405a34910057439100", 878=>X"5d3591006945910000439100003c9140", 879=>X"00459100003c9140733c910000359140", 
    880=>X"6e3c9100003791405f37910069469100", 881=>X"663991006a48910000469100003c9140", 882=>X"57459100004691405946910000489140", 883=>X"00439100003991405c43910000459140", 884=>X"003f91404e3f9100004191405b419100", 
    885=>X"003c9140513c9100003e91404a3e9100", 886=>X"5e489100004a9140503a9100564a9100", 887=>X"004691405c469100003a910000489140", 888=>X"00439140594391000045914060459100", 889=>X"0040914050409100004191404e419100", 
    890=>X"4f3c91005a4c9100003e9140513e9100", 891=>X"003c9100004a91405b4a9100004c9140", 892=>X"004691405c4691000048914056489100", 893=>X"004391404e439100004591405d459100", 894=>X"004091404f409100004191404d419100", 
    895=>X"5d4c9100004d91404a3e91005b4d9100", 896=>X"004a91405c4a9100003e9100004c9140", 897=>X"00469140584691000048914058489100", 898=>X"0043914049439100004591404b459100", 899=>X"4f4091005b4f9100004191404c419100", 
    900=>X"00409100004d9140594d9100004f9140", 901=>X"004a9140594a9100004c9140604c9100", 902=>X"0046914046469100004891405b489100", 903=>X"004391404a4391000045914052459100", 904=>X"4f4d9100005191404b41910058519100", 
    905=>X"004c9140594c910000419100004d9140", 906=>X"4848910055489100004d9140634d9100", 907=>X"00489100004d91406e4d910000489140", 908=>X"004d9140684d9100004c91405e4c9100", 909=>X"594d910000519140494191006d519100", 
    910=>X"004c91405b4c910000419100004d9140", 911=>X"4d48910059489100004d9140694d9100", 912=>X"00489100004d91406f4d910000489140", 913=>X"004d9140674d9100004c91405b4c9100", 914=>X"584c9100004f9140484091006b4f9100", 
    915=>X"004a9140594a910000409100004c9140", 916=>X"4b48910059489100004c9140664c9100", 917=>X"00489100004c9140704c910000489140", 918=>X"004c9140664c9100004a9140634a9100", 919=>X"594c9100004f9140484091006d4f9100", 
    920=>X"004a91405d4a910000409100004c9140", 921=>X"4f4891005a489100004c9140674c9100", 922=>X"00489100004c91406d4c910000489140", 923=>X"004c9140684c9100004a91405f4a9100", 924=>X"414d9100005191403e4191004e519100", 
    925=>X"004c9140434c910000419100004d9140", 926=>X"3e4891003e489100004d9140494d9100", 927=>X"00489100004d91404c4d910000489140", 928=>X"004d91404a4d9100004c9140444c9100", 929=>X"3e4d910000519140404191004f519100", 
    930=>X"004c9140434c910000419100004d9140", 931=>X"404891003f489100004d9140494d9100", 932=>X"00489100004d91404e4d910000489140", 933=>X"004d91404c4d9100004c9140464c9100", 934=>X"424c9100004f91403e4091004b4f9100", 
    935=>X"004a9140414a910000409100004c9140", 936=>X"4148910042489100004c9140424c9100", 937=>X"00489100004c91404a4c910000489140", 938=>X"004c91404c4c9100004a9140414a9100", 939=>X"414c9100004f91403f409100494f9100", 
    940=>X"004a91403d4a910000409100004c9140", 941=>X"414891003d489100004c91404a4c9100", 942=>X"00489100004c91404f4c910000489140", 943=>X"004c9140464c9100004a9140454a9100", 944=>X"694f9100004d91405d3e9100674d9100", 
    945=>X"004d91405d4d9100003e9100004f9140", 946=>X"004a91405a4a9100004c91405a4c9100", 947=>X"004791405b479100004891405a489100", 948=>X"0047914063479100004591405a459100", 949=>X"004791406a479100004391405e439100", 
    950=>X"004d91405b4d9100004a91406d4a9100", 951=>X"004d91405c4d91000051914069519100", 952=>X"0047914057479100004a9140564a9100", 953=>X"00479140664791000043914058439100", 954=>X"004d9140564d9100004a9140684a9100", 
    955=>X"004d9140594d9100005191406b519100", 956=>X"0046914056469100004a91405a4a9100", 957=>X"00469140694691000043914059439100", 958=>X"004c9140584c91000048914069489100", 959=>X"004c9140604c9100004f9140694f9100", 
    960=>X"004691405a4691000048914056489100", 961=>X"004691406e4691000043914058439100", 962=>X"004c9140564c9100004891406a489100", 963=>X"004c91405f4c9100004f9140644f9100", 964=>X"00459140564591000048914051489100", 
    965=>X"004591406d4591000041914052419100", 966=>X"004a91405c4a9100004891406b489100", 967=>X"004a9140584a9100004d91406b4d9100", 968=>X"00459140414591000046914055469100", 969=>X"0045914050459100004191403e419100", 
    970=>X"004a91403c4a9100004691404c469100", 971=>X"004a91403f4a9100004d9140504d9100", 972=>X"004391403d4391000046914041469100", 973=>X"0043914049439100004091403f409100", 974=>X"00499140424991000046914052469100", 
    975=>X"0049914041499100004c91404a4c9100", 976=>X"004391403e439100004691403f469100", 977=>X"00439140504391000040914040409100", 978=>X"004991403e499100004691404c469100", 979=>X"004991403f499100004c91404a4c9100", 
    980=>X"3e519140424591000046914042469100", 981=>X"50499100434f91000045910000519140", 982=>X"00499100005191404f519100004f9140", 983=>X"4f519100004d91404a4a9100404d9100", 984=>X"3b4391003d4c9100004a910000519140", 
    985=>X"00439100005191404c519100004c9140", 986=>X"54519100004a91403c419100394a9100", 987=>X"4f4591003a4991000041910000519140", 988=>X"00459100005191405251910000499140", 989=>X"55519100004a91404a4791003d4a9100", 
    990=>X"48499100404c91000047910000519140", 991=>X"00499100005191404d519100004c9140", 992=>X"4e519100004d91404a4a9100414d9100", 993=>X"4449910032459100004a910000519140", 994=>X"00499100005191405a51910000459140", 
    995=>X"5151910000479140494a910039479100", 996=>X"4f4c91003d499100004a910000519140", 997=>X"004c9100005191405151910000499140", 998=>X"53519100004a9140524d91003d4a9100", 999=>X"424c91003a499100004d910000519140", 
    1000=>X"004c9100005191405451910000499140", 1001=>X"004591403e4591403b4a9100474d9100", 1002=>X"494c91003e499100004d9100004a9100", 1003=>X"004591404b4591000043914044439100", 1004=>X"3e4291403c4a910000499100004c9100", 
    1005=>X"4448910044459100004a910000429140", 1006=>X"004291404a4291000040914041409100", 1007=>X"3d4391003f4691000045910000489100", 1008=>X"0046910000439100003e91403b3e9140", 1009=>X"003c91403f3c91003c42910044459100", 
    1010=>X"0045910000429100003e91404a3e9100", 1011=>X"003a91404b3a91003c43910046469100", 1012=>X"003c9140493c91004045910000469100", 1013=>X"433a9100434391000043910000459100", 1014=>X"423991003c41910000439100003a9140", 
    1015=>X"43379100424091000041910000399140", 1016=>X"43359100423e91000040910000379140", 1017=>X"42349100483d9100003e910000359140", 1018=>X"44329100453b9100003d910000349140", 1019=>X"4531910040399100003b910000329140", 
    1020=>X"002d9140412d91000039910000319140", 1021=>X"003491404d3491000031914049319100", 1022=>X"003a91404b3a9100003791403a379100", 1023=>X"00349140443491000037914043379100", 1024=>X"002d9140442d91000031914040319100", 
    1025=>X"003491404d3491000031914048319100", 1026=>X"003a9140473a91000037914043379100", 1027=>X"00349140463491000037914048379100", 1028=>X"002d9140442d9100003291403d329100", 1029=>X"0035914049359100003291404d329100", 
    1030=>X"003e91404f3e91000039914041399100", 1031=>X"00359140423591000039914043399100", 1032=>X"002d9140402d9100003291403f329100", 1033=>X"0035914049359100003291404a329100", 1034=>X"003e91404e3e9100003991403f399100", 
    1035=>X"00359140443591000039914043399100", 1036=>X"002d91403e2d9100003191403f319100", 1037=>X"003491404b349100003191404d319100", 1038=>X"003a9140463a9100003791403d379100", 1039=>X"00349140433491000037914044379100", 
    1040=>X"002d9140432d91000031914044319100", 1041=>X"003491404e349100003191404b319100", 1042=>X"003a9140483a9100003791403c379100", 1043=>X"00349140433491000037914044379100", 1044=>X"002d9140402d9100003291403e329100", 
    1045=>X"003591404b359100003291404a329100", 1046=>X"003e9140533e91000039914042399100", 1047=>X"00359140433591000039914042399100", 1048=>X"002d9140412d91000032914042329100", 1049=>X"003591404e3591000032914048329100", 
    1050=>X"003e91404f3e91000039914041399100", 1051=>X"00359140423591000039914041399100", 1052=>X"00319140413191000034914040349100", 1053=>X"003791404d3791000034914047349100", 1054=>X"003d91404c3d9100003a91403f3a9100", 
    1055=>X"0037914042379100003a9140473a9100", 1056=>X"00319140433191000034914041349100", 1057=>X"003791404a3791000034914043349100", 1058=>X"003d9140503d9100003a91403e3a9100", 1059=>X"0037914044379100003a9140413a9100", 
    1060=>X"003291403e329100003591403f359100", 1061=>X"003991404d3991000035914049359100", 1062=>X"0041914049419100003e9140433e9100", 1063=>X"0039914043399100003e9140413e9100", 1064=>X"00329140443291000035914043359100", 
    1065=>X"0039914048399100003591404a359100", 1066=>X"004191404f419100003e9140403e9100", 1067=>X"0039914041399100003e9140403e9100", 1068=>X"00319140443191000034914041349100", 1069=>X"0037914046379100003491404c349100", 
    1070=>X"003d9140483d9100003a91403e3a9100", 1071=>X"0037914041379100003a9140473a9100", 1072=>X"00319140413191000034914041349100", 1073=>X"003791404c3791000034914048349100", 1074=>X"003d9140483d9100003a91403b3a9100", 
    1075=>X"0037914041379100003a9140443a9100", 1076=>X"00329140453291000035914041359100", 1077=>X"003991404c399100003591404d359100", 1078=>X"0041914050419100003e9140403e9100", 1079=>X"003991403f399100003e9140423e9100", 
    1080=>X"003291403e3291000035914040359100", 1081=>X"00399140493991000035914049359100", 1082=>X"004191404c419100003e9140433e9100", 1083=>X"0039914040399100003e9140423e9100", 1084=>X"0034914043349100003791403d379100", 
    1085=>X"003a9140493a91000037914045379100", 1086=>X"0040914048409100003d9140403d9100", 1087=>X"003a9140423a9100003d9140423d9100", 1088=>X"00349140433491000037914043379100", 1089=>X"003a9140483a9100003791404a379100", 
    1090=>X"004091404d409100003d9140403d9100", 1091=>X"003a9140443a9100003d9140413d9100", 1092=>X"0035914046359100003991403c399100", 1093=>X"003d9140523d91000039914045399100", 1094=>X"0041914048419100003e9140403e9100", 
    1095=>X"003991403e399100003e9140453e9100", 1096=>X"003e9140423e9100003a9140413a9100", 1097=>X"003791403f379100003a9140433a9100", 1098=>X"00399140403991000035914045359100", 1099=>X"003291403e3291000035914043359100", 
    1100=>X"003291403d329100002d9140412d9100", 1101=>X"002991403f299100002d9140402d9100", 1102=>X"00329140413291000026914045269100", 1103=>X"002f9140472f91000031914043319100", 1104=>X"003a91403d3a91000031914042319100", 
    1105=>X"00379140423791000039914042399100", 1106=>X"00379140423791000035914044359100", 1107=>X"00349140433491000035914043359100", 1108=>X"003a9140403a91000032914040329100", 1109=>X"00379140423791000039914045399100", 
    1110=>X"00379140443791000035914044359100", 1111=>X"00349140473491000035914046359100", 1112=>X"00349120433491000032914045329100", 1113=>X"003791204a3791000035912046359100", 1114=>X"003b9120473b9100003991204b399100", 
    1115=>X"003e91404d3e9100003d9120483d9100", 1116=>X"0040914044409100004191403f419100", 1117=>X"3f39910051459100003e9140403e9100", 1118=>X"003b9120463b91000045910000399140", 1119=>X"003e91204d3e9100003d91204b3d9100", 
    1120=>X"004191204c419100004091204e409100", 1121=>X"004591404d4591000043912047439100", 1122=>X"004c910000439140414391003d4c9100", 1123=>X"004a91000041914047419100444a9100", 1124=>X"00499100004091404040910043499100", 
    1125=>X"494b9100004a91404b4191004e4a9100", 1126=>X"004a910000419120414a9100004b9120", 1127=>X"004691203e4691000048912044489100", 1128=>X"004391203e4391000045912043459100", 1129=>X"00429100003f9140423f914043429100", 
    1130=>X"433c9100003e9140403e910048459100", 1131=>X"46379100003a9140413a9100003c9140", 1132=>X"44439100443b91000045910000379140", 1133=>X"00379140473791000035914041359100", 1134=>X"56489100563c9100003b910000439100", 
    1135=>X"00379140443791000033914043339100", 1136=>X"4047910040439100003c910000489100", 1137=>X"00379140463791000032914043329100", 1138=>X"3f309100504b91000043910000479100", 1139=>X"004b9100003791404b37910000309140", 
    1140=>X"49379100002f9140432f9100404a9100", 1141=>X"3f3091004d4b9100004a910000379140", 1142=>X"004b9100003791404c37910000309140", 1143=>X"4a379100003291404632910042479100", 1144=>X"41339100494891000047910000379140", 
    1145=>X"00489100003791404937910000339140", 1146=>X"4c379100002b91403f2b91003f479100", 1147=>X"432d9100484891000047910000379140", 1148=>X"004891000037914051379100002d9140", 1149=>X"4c379100002f9140422f91004a4a9100", 
    1150=>X"433091004b4b9100004a910000379140", 1151=>X"004b9100003791404f37910000309140", 1152=>X"4a379100002f9140442f9100424a9100", 1153=>X"413091004a4b9100004a910000379140", 1154=>X"004b9100003791404f37910000309140", 
    1155=>X"4b37910000329140463291004a4d9100", 1156=>X"494f910049439100004d910000379140", 1157=>X"3243910000439100004f914041339100", 1158=>X"443291003d4191000043910000339140", 1159=>X"00439100003291404a43910000419140", 
    1160=>X"52439100003f9140483091003f3f9100", 1161=>X"412f91003c3e91000043910000309140", 1162=>X"00439100002f914050439100003e9140", 1163=>X"4f439100003c91404b309100383c9100", 1164=>X"4d3291003f3b91000043910000309140", 
    1165=>X"004391000032914056439100003b9140", 1166=>X"51439100003c9140483391003f3c9100", 1167=>X"483591003e3e91000043910000339140", 1168=>X"004391000035914054439100003e9140", 1169=>X"4c439100003f9140493791003e3f9100", 
    1170=>X"3d2f91003e3791000043910000379140", 1171=>X"00439100002f91405e43910000379140", 1172=>X"54439100003991404630910046399100", 1173=>X"4b329100413b91000043910000309140", 1174=>X"004391000032914052439100003b9140", 
    1175=>X"52439100003c914049339100403c9100", 1176=>X"42329100443b91000043910000339140", 1177=>X"004391000032914052439100003b9140", 1178=>X"57439100003c9140483391003b3c9100", 1179=>X"4a3591003b3e91000043910000339140", 
    1180=>X"004391000035914052439100003e9140", 1181=>X"004f9140583f9100583791005d4f9100", 1182=>X"004f910000379100003f91404c4f9100", 1183=>X"4c4f9100004d9140422f9100454d9100", 1184=>X"434b910043439100004f9100002f9140", 
    1185=>X"4b44910000439100004b914046309100", 1186=>X"00449100004d9100003091404b4d9100", 1187=>X"004a914049329100434a910043419100", 1188=>X"003291404e4b91004e43910000419100", 1189=>X"44489100443f910000439100004b9100", 
    1190=>X"4a4d9100003f9100004891404a339100", 1191=>X"434b910043489100004d910000339140", 1192=>X"484d910000489100004b91403f2d9100", 1193=>X"3d4a91003d419100004d9100002d9140", 1194=>X"5043910000419100004a9140442e9100", 
    1195=>X"00439100004b9100002e9140504b9100", 1196=>X"004891404c3091003d4891003d3f9100", 1197=>X"003091404c4a91004c419100003f9100", 1198=>X"3e4691003e3e910000419100004a9100", 1199=>X"4f4b9100003e91000046914046329100", 
    1200=>X"454a910045469100004b910000329140", 1201=>X"484b910000469100004a91403e2b9100", 1202=>X"47489100473f9100004b9100002b9140", 1203=>X"49419100003f910000489140462d9100", 1204=>X"00419100004a9100002d9140494a9100", 
    1205=>X"00469140472e91003d4691003d3e9100", 1206=>X"002e91404b4891004b3f9100003e9100", 1207=>X"3b4591003b3c9100003f910000489100", 1208=>X"4e4a9100003c9100004591404a309100", 1209=>X"4348910043429100004a910000309140", 
    1210=>X"4a4a9100004291000048914042329100", 1211=>X"4246910042439100004a910000329140", 1212=>X"4845910000439100004691404b379100", 1213=>X"00459100004891000037914048489100", 1214=>X"00459140443291004245910042419100", 
    1215=>X"003291404b4691004b43910000419100", 1216=>X"41439100413f91000043910000469100", 1217=>X"4d439100003f91000043914043339100", 1218=>X"0043910000469100003391404d469100", 1219=>X"00459140432e91004645910046429100", 
    1220=>X"002e91404b4691004b43910000429100", 1221=>X"50489100504591000043910000469100", 1222=>X"414391000045910000489140442d9100", 1223=>X"0043910000469100002d914041469100", 1224=>X"004591404b3091004345910043429100", 
    1225=>X"00309140404391004040910000429100", 1226=>X"413e9140434291000040910000439100", 1227=>X"3d3c91004e45910000429100003e9140", 1228=>X"00459100003e91404b3e9100003c9140", 1229=>X"004a9100003a9140423a9100534a9100", 
    1230=>X"00439100003e91404b3e91003a439100", 1231=>X"00489100003991404139910050489100", 1232=>X"00429100003e91404e3e91003d429100", 1233=>X"0046910000379140463791004e469100", 1234=>X"00439100003e9140513e910042439100", 
    1235=>X"004a91000036914040369100534a9100", 1236=>X"00459100003e9140553e910041459100", 1237=>X"00469100003791404237910047469100", 1238=>X"00439100003e9140513e910044439100", 1239=>X"00459100003991404639910046459100", 
    1240=>X"00429100003e9140523e91003f429100", 1241=>X"00439100003a9140403a91004d439100", 1242=>X"004a9100003e91404b3e9100514a9100", 1243=>X"00429100003291403f32910038429100", 1244=>X"004a9100003e9140593e9100514a9100", 
    1245=>X"00439100003491403f3491003e439100", 1246=>X"004a9100003e9140563e91004f4a9100", 1247=>X"00459100003691404236910042459100", 1248=>X"004a9100003e9140513e91004b4a9100", 1249=>X"0046910000379140443791003c469100", 
    1250=>X"00439100003e9140533e91003d439100", 1251=>X"004a91000036914043369100544a9100", 1252=>X"00459100003e9140513e91003e459100", 1253=>X"00469100003791404537910048469100", 1254=>X"00439100003e9140533e910042439100", 
    1255=>X"00489100003991404139910051489100", 1256=>X"00459100003e91404f3e91003f459100", 1257=>X"44489100004a9140453a91004e4a9100", 1258=>X"463991004a46910000489100003a9140", 1259=>X"00459100003991404645910000469140", 
    1260=>X"00469140413791004337910047469100", 1261=>X"48469100004591000037914046459100", 1262=>X"002b914042439100004691403e2b9100", 1263=>X"00459140473091004945910000439100", 1264=>X"4c489100004691000030914046469100", 
    1265=>X"002d91404e4a910000489140422d9100", 1266=>X"4d3291004a4b9100004a910000379100", 1267=>X"00329140434a9100004b914047369100", 1268=>X"004891403d26910043489100004a9100", 1269=>X"004a91000036910000269140494a9100", 
    1270=>X"004691403e2b91004f3791003e469100", 1271=>X"4845910000489100003791404a489100", 1272=>X"003991404a469100004591404e399100", 1273=>X"003a91404c3a91004543910000469100", 1274=>X"00439100002b91000039914043399100", 
    1275=>X"00379140452b9100473791004f479100", 1276=>X"00479100002b91000035914045359100", 1277=>X"004891404c309100463391004c489100", 1278=>X"4b4d9100004b9100003391404c4b9100", 1279=>X"003f9140474f9100004d91405c3f9100", 
    1280=>X"005091404a3e91004d509100004f9100", 1281=>X"424d9100004f910000309140484f9100", 1282=>X"002f91404d4f9100004d9140442f9100", 1283=>X"453091003e4b9100004f9100003e9100", 1284=>X"003c9140514d9100004b9140453c9100", 
    1285=>X"4b3e9100424a9100004d910000309100", 1286=>X"004b9100003e91404d4b9100004a9140", 1287=>X"49419100003f91404e3f910041489100", 1288=>X"413e91003f4691000048910000419140", 1289=>X"00469100003f91404c3f9100003e9140", 
    1290=>X"4b3f9100003c9140473c910042459100", 1291=>X"423e91004946910000459100003f9140", 1292=>X"4e4391000041914051419100003e9140", 1293=>X"00469100004191404541910000439140", 1294=>X"49419100003f9140403f910041459100", 
    1295=>X"433a9100003e9140433e910000419140", 1296=>X"503f91003f43910000459100003a9140", 1297=>X"443d9100003e91404a3e9100003f9140", 1298=>X"004391000039914042399100003d9140", 1299=>X"463c9100003d91404f3d910046429100", 
    1300=>X"443b91004341910000429100003c9140", 1301=>X"004191000037914042379100003b9140", 1302=>X"453a9100003c9140523c9100423f9100", 1303=>X"433591000039914044399100003a9140", 1304=>X"4a3a9100413e9100003f910000359140", 
    1305=>X"4e3d910051469100003e9100003a9140", 1306=>X"443c91004545910000469100003d9140", 1307=>X"493e91004946910000459100003c9140", 1308=>X"403c91004245910000469100003e9140", 1309=>X"3a3a91004243910000459100003c9140", 
    1310=>X"433991004342910000439100003a9140", 1311=>X"4d3c9100524b91000042910000399140", 1312=>X"413a91004a4a9100004b9100003c9140", 1313=>X"4939910040489100004a9100003a9140", 1314=>X"40379100414691000048910000399140", 
    1315=>X"513c9100555191000046910000379140", 1316=>X"483a9100454f910000519100003c9140", 1317=>X"433991003f4e9100004f9100003a9140", 1318=>X"483a91004d4f9100004e910000399140", 1319=>X"453a9100003c91404b3c9100003a9140", 
    1320=>X"47399100414d9100004f9100003a9140", 1321=>X"4d379100454b9100004d910000399140", 1322=>X"49399100504d9100004b910000379140", 1323=>X"43359100434a9100004d910000399140", 1324=>X"473791004b4b9100004a910000359140", 
    1325=>X"4334910043499100004b910000379140", 1326=>X"0045914041459100004691403f469140", 1327=>X"00499100004391000034914040439100", 1328=>X"423f9140483691004a459100484a9100", 1329=>X"403c9100003e9140423e9100003f9140", 
    1330=>X"004a91000045910000369100003c9140", 1331=>X"413291004a3e91003f42910041489100", 1332=>X"3f3a9100003c9140433c9100003e9140", 1333=>X"003291000039914048399100003a9140", 1334=>X"4a439100484691000048910000429100", 
    1335=>X"48419100004391404f37910047379100", 1336=>X"463e9100003f9140413f910000419140", 1337=>X"00469100003e91000037910000379140", 1338=>X"003991404b399100453d91003f459100", 1339=>X"00459100003d9100003a9140493a9100", 
    1340=>X"00399140443991004b40910050499100", 1341=>X"00499100004091000037914042379100", 1342=>X"00359140423591004a419100494a9100", 1343=>X"004a9100004191000037914048379100", 1344=>X"00349140443491004b439100474c9100", 
    1345=>X"004c910000439100003991404e399100", 1346=>X"0045914042329100494591004b4d9100", 1347=>X"404a91004b4591000043914044439100", 1348=>X"00419100003291403e41910000459140", 1349=>X"004391404c439100414c9100004d9100", 
    1350=>X"0043914044439100004591404b459100", 1351=>X"48469100004a91000045914047459100", 1352=>X"00459140434591000046914046499100", 1353=>X"00459140484591000043914041439100", 1354=>X"3f4191003c459100004c910000499100", 
    1355=>X"484691000045910000419140474a9100", 1356=>X"4343910000469100004391404b439100", 1357=>X"4a459100004391000040914042409100", 1358=>X"3b41910000459100004191404a419100", 1359=>X"003c9140423c9100003e91403d3e9100", 
    1360=>X"4d4d91004c459100004a910000419100", 1361=>X"003991403e399100003a91403c3a9100", 1362=>X"41439100554f910000459100004d9100", 1363=>X"0039914043399100003a91404b3a9100", 1364=>X"494591003e4a9100004f910000439100", 
    1365=>X"00359140473591000037914043379100", 1366=>X"3e43910042499100004a910000459100", 1367=>X"00359140463591000034914043349100", 1368=>X"43419100494a91000049910000439100", 1369=>X"00329140413291000034914043349100", 
    1370=>X"4b4391004a4c9100004a910000419100", 1371=>X"002d9140442d91000031914048319100", 1372=>X"3f419100444a9100004c910000439100", 1373=>X"002d9140432d9100003291404e329100", 1374=>X"3e40910041499100004a910000419100", 
    1375=>X"002d9140412d9100003491404a349100", 1376=>X"4f459100494a91000049910000409100", 1377=>X"002d9140412d91000035914051359100", 1378=>X"4f4691004f4c9100004a910000459100", 1379=>X"002d9140422d9100003791404d379100", 
    1380=>X"44459100464a9100004c910000469100", 1381=>X"002d91403d2d9100003591404e359100", 1382=>X"4443910042499100004a910000459100", 1383=>X"002d91403e2d9100003491404a349100", 1384=>X"41419100474a91000049910000439100", 
    1385=>X"002d9140442d9100003291404d329100", 1386=>X"4d4391004c4c9100004a910000419100", 1387=>X"003991404b3991000031914049319100", 1388=>X"564c91004f4f9100004c910000439100", 1389=>X"0039914050399100002d9140442d9100", 
    1390=>X"484a9100454d9100004f9100004c9100", 1391=>X"00399140513991000032914044329100", 1392=>X"3d459100434a9100004d9100004a9100", 1393=>X"003e9140583e91000035914042359100", 1394=>X"414391003e469100004a910000459100", 
    1395=>X"003e9140573e91000037914047379100", 1396=>X"48439100514c91000046910000439100", 1397=>X"003d9140583d91000034914040349100", 1398=>X"4b459100494a9100004c910000439100", 1399=>X"003e9140593e9100003591403f359100", 
    1400=>X"40419100414a9100004a910000459100", 1401=>X"003e91405f3e9100003291403f329100", 1402=>X"4340910048499100004a910000419100", 1403=>X"004591404e4591000040914045399100", 1404=>X"004591404b4591000043914043439100", 
    1405=>X"004191403e4191004a4a910000499100", 1406=>X"4b4c9100004a9100004591404f459100", 1407=>X"004591404f459100004091403c409100", 1408=>X"003e91403b3e9100494d9100004c9100", 1409=>X"414c9100004d9100004591404e459100", 
    1410=>X"0045914052459100003d91403f3d9100", 1411=>X"003e91403b3e91004d4d9100004c9100", 1412=>X"3b499100004d91000045914050459100", 1413=>X"004591404e459100004091403d409100", 1414=>X"004191403e4191004a4a910000499100", 
    1415=>X"42499100004a9100004591404c459100", 1416=>X"004591405b459100003991403e399100", 1417=>X"003b9140413b91004a4a910000499100", 1418=>X"4b4c9100004a91000045914057459100", 1419=>X"0045914059459100003d9140393d9100", 
    1420=>X"003e91403b3e91004a4d9100004c9100", 1421=>X"454c9100004d91000045914054459100", 1422=>X"0045914051459100003d91403a3d9100", 1423=>X"003e91403e3e9100484d9100004c9100", 1424=>X"4c4f9100004d91000045914051459100", 
    1425=>X"004591404e4591000040914041409100", 1426=>X"005191403e4191004c519100004f9100", 1427=>X"404f910000419100005291404b529100", 1428=>X"005191404c519100004f914045409100", 1429=>X"004d9140443e9100414d910000409100", 
    1430=>X"404c9100003e9100004f9140484f9100", 1431=>X"004d91404e4d9100004c914050439100", 1432=>X"004a914042419100404a910000439100", 1433=>X"4949910000419100004591403b459100", 1434=>X"004591403d4591000049914048409100", 
    1435=>X"004a914046419100504a910000409100", 1436=>X"524c910000419100004591403f459100", 1437=>X"004591403a459100004c91403b3d9100", 1438=>X"004d9140443e9100574d9100003d9100", 1439=>X"504c9100003e9100004591403b459100", 
    1440=>X"004591403d459100004c9140423d9100", 1441=>X"004d9140463e9100524d9100003d9100", 1442=>X"554f9100003e9100004591403c459100", 1443=>X"004591403d459100004f9140423b9100", 1444=>X"005191404c3d910055519100003b9100", 
    1445=>X"544c9100003d91000045914037459100", 1446=>X"004591403d459100004c914053439100", 1447=>X"004d914040419100544d910000439100", 1448=>X"584f910000419100004591403a459100", 1449=>X"0045914035459100004f91403f3e9100", 
    1450=>X"00399140413d910053519100003e9100", 1451=>X"00379140463791000039914049399100", 1452=>X"00519100003d91000039914047399100", 1453=>X"003991404b3991000035914040359100", 1454=>X"00399140493991000034914042349100", 
    1455=>X"003991404a3991000032914045329100", 1456=>X"00399140483991000031914040319100", 1457=>X"003991404d3991000032914041329100", 1458=>X"00399140473991000034914041349100", 1459=>X"003991404a3991000035914042359100", 
    1460=>X"0039914048399100002d9140402d9100", 1461=>X"003991404e399100002f9140422f9100", 1462=>X"003991404c3991000031914044319100", 1463=>X"003991404b3991000032914041329100", 1464=>X"003991404d3991000031914043319100", 
    1465=>X"003991404c3991000032914041329100", 1466=>X"003991404b3991000034914043349100", 1467=>X"564391003e4c91000035914042359100", 1468=>X"48419100434a9100004c910000439140", 1469=>X"444091003f499100004a910000419140", 
    1470=>X"4e4191004e4a91000049910000409140", 1471=>X"004a9100003d9140403d910000419140", 1472=>X"003591403c4d9140423591004f3e9100", 1473=>X"004c914045379100424c9100004d9100", 1474=>X"4d4f9100004d910000379140494d9100", 
    1475=>X"003491404f519100004f914044349100", 1476=>X"423d91004552910000519100003e9100", 1477=>X"0039914044519100005291404e399100", 1478=>X"004f91403c2d9100454f910000519100", 1479=>X"00519100003d9100002d914049519100", 
    1480=>X"003e91404b329100443e9100444d9100", 1481=>X"414c9100004d91000045914050459100", 1482=>X"0032914049499100004791404f479100", 1483=>X"4d4a9100424a9100004c910000499100", 1484=>X"004a9100004c9140464c9100004a9140", 
    1485=>X"004d9140402d910042489100444d9100", 1486=>X"00489100004b9100002d9140444b9100", 1487=>X"004a9140492e910036419100434a9100", 1488=>X"4646910000489100002e914041489100", 1489=>X"002b91404445910000469140442b9100", 
    1490=>X"004391404d3091003f43910000459100", 1491=>X"00419100004591000030914047459100", 1492=>X"004691403c2491003d3f91004e469100", 1493=>X"4145910000489100002491404d489100", 1494=>X"003c9140403c9100003f91404a299100", 
    1495=>X"00299140423591000039914041399100", 1496=>X"00399140443991000045910000359100", 1497=>X"4b3f91003d489100003c91404b3c9100", 1498=>X"002d9140463c9100003f9140422d9100", 1499=>X"003e9140422e91004e3e9100003c9100", 
    1500=>X"4646910000489100003a9140433a9100", 1501=>X"002e91403e3291000037914041379100", 1502=>X"003791404b3791000046910000329100", 1503=>X"4f3e9100414f9100003a9140443a9100", 1504=>X"002e914051439100003e9140392e9100", 
    1505=>X"564891003b4b9100004f910000439100", 1506=>X"464d9100004b91000048914043309100", 1507=>X"404a9100004d9100004a91404e4a9100", 1508=>X"4a4b9100004a9100004691403f469100", 1509=>X"004b9100004891000030914049489100", 
    1510=>X"00489100004591404045910044489100", 1511=>X"00469100004391404643910043469100", 1512=>X"00429140412d91004442910044459100", 1513=>X"002d9140394091004143910000459100", 1514=>X"443e9100443691000043910000409100", 
    1515=>X"3f32910000369100003e914040269100", 1516=>X"49379100003691404b36910000329140", 1517=>X"003991403e3991000037910000269140", 1518=>X"0039914043399100003e9140513e9100", 1519=>X"41269100443691000037914046379100", 
    1520=>X"43369100003291404532910000369140", 1521=>X"00379100002691404a37910000369140", 1522=>X"003e91404f3e91000039914040399100", 1523=>X"00369140413691000039914044399100", 1524=>X"40329100003791404026910043379100", 
    1525=>X"49399100003791404b37910000329140", 1526=>X"003a91403f3a91000039910000269140", 1527=>X"003a9140413a9100003e9140503e9100", 1528=>X"3a269100433791000039914045399100", 1529=>X"4e379100003291403f32910000379140", 
    1530=>X"00399100002691404939910000379140", 1531=>X"003e91404b3e9100003a9140443a9100", 1532=>X"003a9140443a9100003c9140443c9100", 1533=>X"44369100003991403e2691003d399100", 1534=>X"483a9100003991404539910000369140", 
    1535=>X"003c91403b3c9100003a910000269140", 1536=>X"003c9140413c9100003f91404b3f9100", 1537=>X"402691003f399100003a9140433a9100", 1538=>X"46399100003691404936910000399140", 1539=>X"003a910000269140473a910000399140", 
    1540=>X"003f91404a3f9100003c91403f3c9100", 1541=>X"003a9140433a9100003c91403f3c9100", 1542=>X"493a9100003991404126910043399100", 1543=>X"4f429100003e91404f3e9100003a9140", 1544=>X"00439140484391000042910000269140", 
    1545=>X"0043914044439100004691404f469100", 1546=>X"3d269100443a9100003e91403a3e9100", 1547=>X"483a91000037914044379100003a9140", 1548=>X"003e9100002691404c3e9100003a9140", 1549=>X"004691404e469100004391404e439100", 
    1550=>X"003e91403c3e91000043914041439100", 1551=>X"42399100003c914042269100403c9100", 1552=>X"4d3f9100003c91404c3c910000399140", 1553=>X"0042914045429100003f910000269140", 1554=>X"004291403e429100004591404a459100", 
    1555=>X"402691003d3c9100003f9140423f9100", 1556=>X"4c3c91000039914047399100003c9140", 1557=>X"003f9100002691404d3f9100003c9140", 1558=>X"004591404a4591000042914043429100", 1559=>X"003f9140403f91000042914041429100", 
    1560=>X"00329140403291403c3e91003c369100", 1561=>X"003091404730910000369100003e9100", 1562=>X"3f439100444a91000032914048329100", 1563=>X"0032914048329100002e9140412e9100", 1564=>X"494291003e489100004a910000439100", 
    1565=>X"4b329100002d91403f2d910049459100", 1566=>X"00489100004291000045910000329140", 1567=>X"002b9140402b91004043910040469100", 1568=>X"00359140423591000037914051379100", 1569=>X"0046910000439100003791404b379100", 
    1570=>X"4633910044439100443f91004e489100", 1571=>X"00439100003791404e37910000339140", 1572=>X"4f479100484a910000489100003f9100", 1573=>X"003791404c3791000032914046329100", 1574=>X"4d4391004c4b9100004a910000479100", 
    1575=>X"4530910000309140423091004d489100", 1576=>X"49309100002e9140482e910000309140", 1577=>X"004b9100004391000048910000309140", 1578=>X"002d9140462d910045489100464d9100", 1579=>X"004d910000489100003091404b309100", 
    1580=>X"442b9100544c9100544691004d4f9100", 1581=>X"004c9100003091404b309100002b9140", 1582=>X"4d45910049519100004f910000469100", 1583=>X"4d35910000299140422991004d4d9100", 1584=>X"4a359100003391404733910000359140", 
    1585=>X"0051910000459100004d910000359140", 1586=>X"0032914043329100344691003f4d9100", 1587=>X"004d910000469100003591404a359100", 1588=>X"413091004c4891004c4591003f4b9100", 1589=>X"00489100003591404935910000309140", 
    1590=>X"43469100434a9100004b910000459100", 1591=>X"494b910049439100004a9140422e9100", 1592=>X"0046910000439100004b9100002e9140", 1593=>X"004a91404b339100414a910041419100", 1594=>X"003391403f4891003f3f910000419100", 
    1595=>X"3e4691003e3e9100003f910000489100", 1596=>X"4c3f9100003e91000046914049359100", 1597=>X"003f910000489100003591404c489100", 1598=>X"004691403f29910045469100453e9100", 1599=>X"002991403f4591003f3c9100003e9100", 
    1600=>X"41439100413a9100003c910000459100", 1601=>X"533f9100003a910000439140492b9100", 1602=>X"003f910000489100002b914053489100", 1603=>X"004691404b30910045469100453e9100", 1604=>X"0030914042459100423c9100003e9100", 
    1605=>X"42439100423a9100003c910000459100", 1606=>X"4e3c9100003a91000043914049329100", 1607=>X"003c910000459100003291404e459100", 1608=>X"004391403b26910044439100443a9100", 1609=>X"002691404142910041399100003a9100", 
    1610=>X"4b4391004b3a91000039910000429100", 1611=>X"40399100003a910000439140462b9100", 1612=>X"42379100003991000041914040419100", 1613=>X"42359100003791000040914042409100", 1614=>X"00359100003e9100002b9140423e9100", 
    1615=>X"002d9140422d9140433d910043349100", 1616=>X"4d4091004d37910000349100003d9100", 1617=>X"002d9140462d9100002b9140432b9100", 1618=>X"4d4191004d3991000037910000409100", 1619=>X"4c3b910000399100004191403c299100", 
    1620=>X"003b910000439100002991404c439100", 1621=>X"004591404226910049459100493d9100", 1622=>X"002691404b4791004b3e9100003d9100", 1623=>X"4849910048409100003e910000479100", 1624=>X"4741910000409100004991404f2d9100", 
    1625=>X"4c43910000419100004a9140474a9100", 1626=>X"4b45910000439100004c91404c4c9100", 1627=>X"00459100004d9100002d91404b4d9100", 1628=>X"46910081472691003f4691004a4f9100", 1629=>X"45914042459100414d9100004f910000", 
    1630=>X"43914042439100404c9100004d910000", 1631=>X"41914044419100484a9100004c910000", 1632=>X"499100004a9100004591404b45910000", 1633=>X"4591404d459100004091403b40910040", 1634=>X"3e91403c3e9100504a91000049910000", 
    1635=>X"4c9100004a9100004591405045910000", 1636=>X"4591404a459100003d9140393d910048", 1637=>X"3e91403e3e91004a4d9100004c910000", 1638=>X"4f9100004d9100004591405145910000", 1639=>X"4591405145910000409140434091004c", 
    1640=>X"419140434191004f519100004f910000", 1641=>X"49910000519100004591404c45910000", 1642=>X"4591405a459100003991403f39910038", 1643=>X"3b9140403b9100474a91000049910000", 1644=>X"4c9100004a9100004591405245910000", 
    1645=>X"26914054459100003d9140373d91004a", 1646=>X"3e91004a4d9100004c91000045910000", 1647=>X"4d9100004591404d459100003e91403c", 1648=>X"459100003d91403b3d91003d4c910000", 1649=>X"3e91004c4d9100004c91000045914055", 
    1650=>X"4d91000045914050459100003e91403d", 1651=>X"459100003b91403f3b9100434a910000", 1652=>X"4991004a4c9100004a9100004591405a", 1653=>X"910000499100002d910081402d910050", 1654=>X"0081422991003f459100444a9100004c", 
    1655=>X"00454a9100004a910000459100002991", 1656=>X"002b9100814c2b910049469100494391", 1657=>X"41499100004a91000043910000469100", 1658=>X"2d910081432d91004245910042409100", 1659=>X"4a910000499100004091000045910000", 
    1660=>X"91008142299100474591004741910045", 1661=>X"9100004a910000419100004591000029", 1662=>X"0081452691004f4a91004f4591004b4d", 1663=>X"00004d910000459100004a9100002691", 1664=>X"81492b9100464a910046469100444c91", 
    1665=>X"4245910000469100004a9100002b9100", 1666=>X"489100002d9100814d2d910042489100", 1667=>X"4191003c4a9100004c91000045910000", 1668=>X"ff40834b3591004b2e91005a3e910039", 1669=>X"00359140404b4c0351ff00404b4c0351", 
    1670=>X"004a910000419100003e9100002e9100", 1671=>X"912036140d0351ff0036140d0351ff00", 1672=>X"9100004f91204a4f9100004d9120404d", 1673=>X"9100005291204b529100005191204f51", 1674=>X"91000046912048469100004591203e45", 
    1675=>X"9100004a9120504a9100004891204a48", 1676=>X"9100004a91204a4a9100004891204048", 1677=>X"9100004d91204c4d9100004b9120484b", 1678=>X"91000043912048439100004191203a41", 1679=>X"91000046912046469100004591204a45", 
    1680=>X"9100004691204a469100004591204045", 1681=>X"9100004a91204b4a9100004891204e48", 1682=>X"91000043912040439100004591203f45", 1683=>X"9100003f9120443f9100004191204541", 1684=>X"9100004591204f459100004391204443", 
    1685=>X"91000048912054489100004691204a46", 1686=>X"91000041912042419100004391203f43", 1687=>X"9100003e9120423e9100003f9120423f", 1688=>X"9100004391204b439100004191203a41", 1689=>X"91000046912046469100004591204a45", 
    1690=>X"9100003a9120443a9100003991204339", 1691=>X"9100003e91204a3e9100003c91204f3c", 1692=>X"9100003e91204b3e9100003c91203f3c", 1693=>X"9100004191204c419100003f91204c3f", 1694=>X"91000037912047379100003591204135", 
    1695=>X"9100003a91203e3a9100003991204839", 1696=>X"9100003a9120483a9100003991203f39", 1697=>X"9100003e91204d3e9100003c9120483c", 1698=>X"9100003a9120413a9100003c91203d3c", 1699=>X"91000037912044379100003991204239", 
    1700=>X"9100003c91204b3c9100003a91203c3a", 1701=>X"9100003f91204c3f9100003e9120493e", 1702=>X"9100003c91203d3c9100003e91203f3e", 1703=>X"91000039912041399100003a9120453a", 1704=>X"9100003e91204e3e9100003c91203d3c", 
    1705=>X"9100004291204d429100004091204940", 1706=>X"9100003e91203e3e9100003f91203c3f", 1707=>X"9100003a9120443a9100003c9120403c", 1708=>X"91000043912049439100004291203e42", 1709=>X"91203f48912043469100004591204d45", 
    1710=>X"9100004a91203d379100484a91000048", 1711=>X"91000046910000439100003791203a43", 1712=>X"91003c4391003c409100544c91005446", 1713=>X"824735910000319100843b3191006c3d", 1714=>X"004c91000040910000439100003d9100", 
    1715=>X"45419100414a91004145910000469100", 1716=>X"9100814332910000359100814d3e9100", 1717=>X"91000045910000419100003e91000032", 1718=>X"9100452c910046419100463e91004647", 1719=>X"0000419100002c9100003b910084453b", 
    1720=>X"403b38914000479100004a9100003e91", 1721=>X"403d359100003b9140483b9100003891", 1722=>X"4044329100003891404d389100003591", 1723=>X"40402f9100003591404c359100003291", 1724=>X"40442c9100003291404a329100002f91", 
    1725=>X"43289100002d910081462d9100002c91", 1726=>X"449100404091003d4a91003d47910081", 1727=>X"91008150389100503491004c3b910040", 1728=>X"910000449100003b9100003491000038", 1729=>X"91004040910000479100004a91000040", 
    1730=>X"9100453491004f3c91004b4591004048", 1731=>X"00004391404143910000459100834539", 1732=>X"00004091000041910000399140404191", 1733=>X"00404b4c0351ff408343379100454091", 1734=>X"91000037910000289140404b4c0351ff", 
    1735=>X"ff000040910000489100003c91000034", 1736=>X"4243912036140d0351ff0036140d0351", 1737=>X"4a439100004191203f41910000439120", 1738=>X"42409100004091204040910000439120", 1739=>X"49409100003e9120443e910000409120", 
    1740=>X"3d459100003c9120433c910000409120", 1741=>X"4d459100004391204043910000459120", 1742=>X"3d419100004191203f41910000459120", 1743=>X"49419100004091204040910000419120", 1744=>X"41479100003e9120433e910000419120", 
    1745=>X"49479100004591204045910000479120", 1746=>X"41439100004391204143910000479120", 1747=>X"48439100004191204441910000439120", 1748=>X"41489100004091204140910000439120", 1749=>X"49489100004791204347910000489120", 
    1750=>X"404a9100004591203b45910000489120", 1751=>X"4a4a91000048912041489100004a9120", 1752=>X"414c91000047912040479100004a9120", 1753=>X"494c9100004a9120474a9100004c9120", 1754=>X"414d9100004891203d489100004c9120", 
    1755=>X"464d9100004c9120444c9100004d9120", 1756=>X"3f4f9100004a9120414a9100004d9120", 1757=>X"4a4f9100004d91203e4d9100004f9120", 1758=>X"3f489100004c9120434c9100004f9120", 1759=>X"4a489100004791203f47910000489120", 
    1760=>X"424a9100004591204145910000489120", 1761=>X"4c4a91000048912040489100004a9120", 1762=>X"3d4491000047912041479100004a9120", 1763=>X"4d449100004291203f42910000449120", 1764=>X"3a489100004091204440910000449120", 
    1765=>X"44489100004791204547910000489120", 1766=>X"44419100004591203d45910000489120", 1767=>X"48419100004091204340910000419120", 1768=>X"3e479100003e9120423e910000419120", 1769=>X"4a479100004591204245910000479120", 
    1770=>X"3c459100003c91203e3c910000479120", 1771=>X"52459100004391203d43910000459120", 1772=>X"40449100003b91203e3b910000459120", 1773=>X"48449100004291203e42910000449120", 1774=>X"403c9100004091204040910000449120", 
    1775=>X"47399100003b91203f3b9100003c9120", 1776=>X"433e9100003891204638910000399120", 1777=>X"473b9100003c9120443c9100003e9120", 1778=>X"41409100003991203f399100003b9120", 1779=>X"433c9100003e9120403e910000409120", 
    1780=>X"3e419100003b9120413b9100003c9120", 1781=>X"433e9100004091204440910000419120", 1782=>X"3e439100003c9120423c9100003e9120", 1783=>X"43409100004191203c41910000439120", 1784=>X"40459100003e91203d3e910000409120", 
    1785=>X"42419100004391203f43910000459120", 1786=>X"3e439100004091203f40910000419120", 1787=>X"4c479100004591204a45910000439120", 1788=>X"4091003f3c9100814748910000479120", 1789=>X"91008141379100413491003f4391003f", 
    1790=>X"91000040910000439100003491000037", 1791=>X"9100494091004b49910000489100003c", 1792=>X"00003991008146399100463791004945", 1793=>X"00004991000040910000459100003791", 1794=>X"00003d91204e3d9100003991203f3991", 
    1795=>X"00004591203d459100004091204d4091", 1796=>X"3f4091004749910000499100814a4991", 1797=>X"399100813e3991003e3791003f459100", 1798=>X"49910000409100004591000037910000", 1799=>X"45910048419100483e91004c4a910000", 
    1800=>X"91000039910081473991004735910048", 1801=>X"9100003e910000419100004591000035", 1802=>X"91204f3e9100003991203f399100004a", 1803=>X"912042459100004191204b419100003e", 1804=>X"00464a9100004a9100814e4a91000045", 
    1805=>X"8140399100403591003e4591003e4191", 1806=>X"00419100004591000035910000399100", 1807=>X"40439100403e910046479100004a9100", 1808=>X"35910000379100814837910048359100", 1809=>X"37910000479100003e91000043910000", 
    1810=>X"3e9100003b91204d3b91000037912044", 1811=>X"479100004391203f439100003e91204c", 1812=>X"9100403e910049479100004791008150", 1813=>X"00003791008145379100453591004043", 1814=>X"0000479100003e910000439100003591", 
    1815=>X"004934910048439100484091004c4891", 1816=>X"00439100003491000037910081493791", 1817=>X"003791203b3791000048910000409100", 1818=>X"004091204d409100003c91204d3c9100", 1819=>X"48910081504891000043912040439100", 
    1820=>X"3491003f4391003f4091004848910000", 1821=>X"91000034910000379100813c3791003c", 1822=>X"91003c45910000489100004091000043", 1823=>X"0081453991004534910041419100413c", 1824=>X"00003c91000041910000349100003991", 
    1825=>X"204d3991000035912042359100004591", 1826=>X"203e419100003c9120503c9100003991", 1827=>X"4845910000459100814d459100004191", 1828=>X"3e3591003e3491003c4191003c3c9100", 1829=>X"3c910000419100003491000035910081", 
    1830=>X"419100453e91004e4691000045910000", 1831=>X"91000035910081453591004532910045", 1832=>X"910000469100003e9100004191000032", 1833=>X"9100003a91204d3a9100003591204635", 1834=>X"9100004191203d419100003e9120503e", 
    1835=>X"00403e91004546910000469100814f46", 1836=>X"00359100814135910041329100404191", 1837=>X"00469100003e91000041910000329100", 1838=>X"45349100453191004b43910047469100", 1839=>X"46910000439100003191000034910081", 
    1840=>X"3791204a379100003491204634910000", 1841=>X"3d9120423d9100003a9120493a910000", 1842=>X"91004b46910000469100815546910000", 1843=>X"91003f3191004143910041409100413d", 1844=>X"00004391000031910000349100813f34", 
    1845=>X"004145910000469100003d9100004091", 1846=>X"81473691004730910049429100493e91", 1847=>X"003e9100004291000030910000369100", 1848=>X"4e399100003291203e32910000459100", 1849=>X"41429100003e91204d3e910000399120", 
    1850=>X"45910000459100814c45910000429120", 1851=>X"369100423091003d4291003d3e91004a", 1852=>X"91000042910000309100003691008142", 1853=>X"9100413791003d3e91003d3a9100003e", 1854=>X"004443910000459100002b9100823e2b", 
    1855=>X"003e910000379100002e9100824d2e91", 1856=>X"4b3a910049409100493d9100003a9100", 1857=>X"409100003a910000289100823c289100", 1858=>X"3e91004141910000439100003d910000", 1859=>X"9100824d299100493991003e3e910042", 
    1860=>X"910000419100003e9100003991000029", 1861=>X"00003e9100824b3991004b2d91003f40", 1862=>X"00409100002d91000039910082453c91", 1863=>X"3591008242359100422e9100413e9100", 1864=>X"2b9100423a9100003c9100002e910000", 
    1865=>X"910047399100003a9100002b9100823d", 1866=>X"ff00404b4c0351ff40874d3591004d26", 1867=>X"3991000026910000359140404b4c0351", 1868=>X"0351ff0040420f0351ff00003e910000", 1869=>X"0351ff0040420f0351002fff0140420f",
    -- End of bach_tocatta_fugue_d_minor.mid

-- OneDividedByDivision Constants
1870=>X"00040000000555550008000000100000", 1871=>X"00020000000249250002aaab00033333", 1872=>X"000155550001745d0001999a0001c71c", 1873=>X"00010000000111110001249200013b14", 1874=>X"0000cccd0000d7940000e38e0000f0f1", 
1875=>X"0000aaab0000b2160000ba2f0000c30c", 1876=>X"00009249000097b400009d8a0000a3d7", 1877=>X"00008000000084210000888900008d3e", 1878=>X"000071c7000075070000787800007c1f", 1879=>X"000066660000690700006bca00006eb4", 
1880=>X"00005d1700005f4100006186000063e7", 1881=>X"00005555000057260000590b00005b06", 1882=>X"00004ec500005050000051ec00005398", 1883=>X"0000492500004a7900004bda00004d48", 1884=>X"000044440000456c0000469f000047dc", 
1885=>X"00004000000041040000421100004326", 1886=>X"00003c3c00003d2200003e1000003f04", 1887=>X"000038e4000039b100003a8400003b5d", 1888=>X"000035e50000369d0000375a0000381c", 1889=>X"00003333000033d90000348300003532", 
1890=>X"000030c300003159000031f400003291", 1891=>X"00002e8c00002f1500002fa100003030", 1892=>X"00002c8600002d0300002d8300002e06", 1893=>X"00002aab00002b1e00002b9300002c0b", 1894=>X"000028f600002960000029cc00002a3a", 
1895=>X"00002762000027c4000028280000288e", 1896=>X"000025ed00002648000026a400002702", 1897=>X"00002492000024e70000253d00002594", 1898=>X"0000234f0000239e000023ee0000243f", 1899=>X"000022220000226c000022b600002302", 
1900=>X"000021080000214d00002193000021da", 1901=>X"000020000000204100002082000020c5", 1902=>X"00001f0800001f4400001f8200001fc0", 1903=>X"00001e1e00001e5700001e9100001ecc", 1904=>X"00001d4200001d7800001dae00001de6", 
1905=>X"00001c7200001ca500001cd800001d0d", 1906=>X"00001bad00001bdd00001c0e00001c40", 1907=>X"00001af300001b2000001b4f00001b7d", 1908=>X"00001a4200001a6d00001a9900001ac5", 1909=>X"0000199a000019c3000019ed00001a17", 
1910=>X"000018fa000019210000194900001971", 1911=>X"0000186200001887000018ad000018d3", 1912=>X"000017d0000017f4000018180000183d", 1913=>X"00001746000017680000178a000017ad", 1914=>X"000016c1000016e20000170300001724", 
1915=>X"000016430000166200001681000016a1", 1916=>X"000015ca000015e70000160600001624", 1917=>X"00001555000015720000158f000015ac", 1918=>X"000014e6000015010000151d00001539", 1919=>X"0000147b00001495000014b0000014cb", 
1920=>X"000014140000142d0000144700001461", 1921=>X"000013b1000013ca000013e2000013fb", 1922=>X"000013520000136a0000138100001399", 1923=>X"000012f70000130d000013240000133b", 1924=>X"0000129e000012b4000012ca000012e0", 
1925=>X"000012490000125e0000127300001289", 1926=>X"000011f70000120b0000122000001234", 1927=>X"000011a8000011bb000011cf000011e3", 1928=>X"0000115b0000116e0000118100001194", 1929=>X"00001111000011230000113600001148", 
1930=>X"000010c9000010db000010ed000010ff", 1931=>X"0000108400001095000010a7000010b8", 1932=>X"00001041000010520000106200001073", 1933=>X"00001000000010100000102000001031", 1934=>X"00000fc100000fd100000fe000000ff0", 
1935=>X"00000f8400000f9300000fa200000fb2", 1936=>X"00000f4900000f5700000f6600000f75", 1937=>X"00000f0f00000f1d00000f2c00000f3a", 1938=>X"00000ed700000ee500000ef300000f01", 1939=>X"00000ea100000eae00000ebc00000ec9", 
1940=>X"00000e6c00000e7900000e8600000e94", 1941=>X"00000e3900000e4600000e5200000e5f", 1942=>X"00000e0700000e1300000e2000000e2c", 1943=>X"00000dd600000de200000def00000dfb", 1944=>X"00000da700000db300000dbf00000dcb", 
1945=>X"00000d7900000d8500000d9000000d9c", 1946=>X"00000d4c00000d5800000d6300000d6e", 1947=>X"00000d2100000d2c00000d3700000d41", 1948=>X"00000cf600000d0100000d0b00000d16", 1949=>X"00000ccd00000cd700000ce100000cec", 
1950=>X"00000ca400000cae00000cb800000cc3", 1951=>X"00000c7d00000c8700000c9000000c9a", 1952=>X"00000c5600000c6000000c6a00000c73", 1953=>X"00000c3100000c3a00000c4300000c4d", 1954=>X"00000c0c00000c1500000c1e00000c28", 
1955=>X"00000be800000bf100000bfa00000c03", 1956=>X"00000bc500000bce00000bd700000bdf", 1957=>X"00000ba300000bab00000bb400000bbd", 1958=>X"00000b8100000b8a00000b9200000b9a", 1959=>X"00000b6100000b6900000b7100000b79", 
1960=>X"00000b4100000b4900000b5100000b59", 1961=>X"00000b2100000b2900000b3100000b39", 1962=>X"00000b0300000b0a00000b1200000b1a", 1963=>X"00000ae500000aec00000af400000afb", 1964=>X"00000ac700000acf00000ad600000add", 
1965=>X"00000aab00000ab200000ab900000ac0", 1966=>X"00000a8f00000a9500000a9d00000aa4", 1967=>X"00000a7300000a7a00000a8100000a88", 1968=>X"00000a5800000a5f00000a6500000a6c", 1969=>X"00000a3d00000a4400000a4b00000a51", 
1970=>X"00000a2300000a2a00000a3000000a37", 1971=>X"00000a0a00000a1000000a1700000a1d", 1972=>X"000009f1000009f7000009fe00000a04", 1973=>X"000009d9000009df000009e5000009eb", 1974=>X"000009c1000009c7000009cd000009d3", 
1975=>X"000009a9000009af000009b5000009bb", 1976=>X"00000992000009980000099d000009a3", 1977=>X"0000097b00000981000009870000098c", 1978=>X"000009650000096b0000097000000976", 1979=>X"0000094f000009550000095a0000095f", 
1980=>X"0000093a0000093f000009440000094a", 1981=>X"000009250000092a0000092f00000934", 1982=>X"00000910000009150000091a0000091f", 1983=>X"000008fc00000901000009060000090b", 1984=>X"000008e8000008ec000008f1000008f6", 
1985=>X"000008d4000008d9000008de000008e3", 1986=>X"000008c1000008c5000008ca000008cf", 1987=>X"000008ae000008b2000008b7000008bc", 1988=>X"0000089b000008a0000008a4000008a9", 1989=>X"000008890000088d0000089200000896", 
1990=>X"000008760000087b0000087f00000884", 1991=>X"00000865000008690000086e00000872", 1992=>X"00000853000008580000085c00000860", 1993=>X"00000842000008460000084b0000084f", 1994=>X"00000831000008350000083a0000083e", 
1995=>X"0000082100000825000008290000082d", 1996=>X"0000081000000814000008180000081c", 1997=>X"0000080000000804000008080000080c", 1998=>X"000007f0000007f4000007f8000007fc", 1999=>X"000007e0000007e4000007e8000007ec", 
2000=>X"000007d1000007d5000007d9000007dd", 2001=>X"000007c2000007c6000007c9000007cd", 2002=>X"000007b3000007b7000007ba000007be", 2003=>X"000007a4000007a8000007ac000007af", 2004=>X"00000796000007990000079d000007a1", 
2005=>X"000007880000078b0000078f00000792", 2006=>X"000007790000077d0000078000000784", 2007=>X"0000076c0000076f0000077300000776", 2008=>X"0000075e000007610000076500000768", 2009=>X"0000075000000754000007570000075b", 
2010=>X"00000743000007460000074a0000074d", 2011=>X"00000736000007390000073d00000740", 2012=>X"000007290000072c0000073000000733", 2013=>X"0000071c000007200000072300000726", 2014=>X"00000710000007130000071600000719", 
2015=>X"00000704000007070000070a0000070d", 2016=>X"000006f7000006fa000006fd00000700", 2017=>X"000006eb000006ee000006f1000006f4", 2018=>X"000006df000006e2000006e5000006e8", 2019=>X"000006d4000006d7000006d9000006dc", 
2020=>X"000006c8000006cb000006ce000006d1", 2021=>X"000006bd000006bf000006c2000006c5", 2022=>X"000006b1000006b4000006b7000006ba", 2023=>X"000006a6000006a9000006ac000006af", 2024=>X"0000069b0000069e000006a1000006a3", 
2025=>X"00000690000006930000069600000699", 2026=>X"00000686000006880000068b0000068e", 2027=>X"0000067b0000067e0000068000000683", 2028=>X"00000671000006730000067600000679", 2029=>X"00000666000006690000066c0000066e", 
2030=>X"0000065c0000065f0000066100000664", 2031=>X"0000065200000655000006570000065a", 2032=>X"000006480000064b0000064d00000650", 2033=>X"0000063e000006410000064300000646", 2034=>X"00000635000006370000063a0000063c", 
2035=>X"0000062b0000062e0000063000000632", 2036=>X"00000622000006240000062600000629", 2037=>X"000006180000061b0000061d0000061f", 2038=>X"0000060f000006110000061400000616", 2039=>X"00000606000006080000060b0000060d", 
2040=>X"000005fd000005ff0000060200000604", 2041=>X"000005f4000005f6000005f9000005fb", 2042=>X"000005eb000005ed000005f0000005f2", 2043=>X"000005e3000005e5000005e7000005e9", 2044=>X"000005da000005dc000005de000005e0", 
2045=>X"000005d1000005d4000005d6000005d8", 2046=>X"000005c9000005cb000005cd000005cf", 2047=>X"000005c1000005c3000005c5000005c7", 2048=>X"000005b8000005bb000005bd000005bf", 2049=>X"000005b0000005b2000005b4000005b6", 
2050=>X"000005a8000005aa000005ac000005ae", 2051=>X"000005a0000005a2000005a4000005a6", 2052=>X"000005980000059a0000059c0000059e", 2053=>X"00000591000005930000059500000597", 2054=>X"000005890000058b0000058d0000058f", 
2055=>X"00000581000005830000058500000587", 2056=>X"0000057a0000057c0000057e0000057f", 2057=>X"00000572000005740000057600000578", 2058=>X"0000056b0000056d0000056f00000571", 2059=>X"00000564000005660000056700000569", 
2060=>X"0000055c0000055e0000056000000562", 2061=>X"0000055500000557000005590000055b", 2062=>X"0000054e000005500000055200000554", 2063=>X"00000547000005490000054b0000054d", 2064=>X"00000540000005420000054400000546", 
2065=>X"000005390000053b0000053d0000053f", 2066=>X"00000533000005340000053600000538", 2067=>X"0000052c0000052e0000052f00000531", 2068=>X"0000052500000527000005290000052a", 2069=>X"0000051f000005200000052200000524", 
2070=>X"000005180000051a0000051b0000051d", 2071=>X"00000512000005130000051500000517", 2072=>X"0000050b0000050d0000050f00000510", 2073=>X"0000050500000507000005080000050a", 2074=>X"000004ff000005000000050200000503", 
2075=>X"000004f9000004fa000004fc000004fd", 2076=>X"000004f2000004f4000004f5000004f7", 2077=>X"000004ec000004ee000004ef000004f1", 2078=>X"000004e6000004e8000004e9000004eb", 2079=>X"000004e0000004e2000004e3000004e5", 
2080=>X"000004da000004dc000004dd000004df", 2081=>X"000004d5000004d6000004d7000004d9", 2082=>X"000004cf000004d0000004d2000004d3", 2083=>X"000004c9000004ca000004cc000004cd", 2084=>X"000004c3000004c5000004c6000004c8", 
2085=>X"000004be000004bf000004c0000004c2", 2086=>X"000004b8000004b9000004bb000004bc", 2087=>X"000004b2000004b4000004b5000004b7", 2088=>X"000004ad000004ae000004b0000004b1", 2089=>X"000004a8000004a9000004aa000004ac", 
2090=>X"000004a2000004a4000004a5000004a6", 2091=>X"0000049d0000049e0000049f000004a1", 2092=>X"00000498000004990000049a0000049c", 2093=>X"00000492000004940000049500000496", 2094=>X"0000048d0000048e0000049000000491", 
2095=>X"00000488000004890000048b0000048c", 2096=>X"00000483000004840000048500000487", 2097=>X"0000047e0000047f0000048000000482", 2098=>X"000004790000047a0000047b0000047c", 2099=>X"00000474000004750000047600000477", 
2100=>X"0000046f000004700000047100000473", 2101=>X"0000046a0000046b0000046c0000046e", 2102=>X"00000465000004660000046800000469", 2103=>X"00000460000004610000046300000464", 2104=>X"0000045c0000045d0000045e0000045f", 
2105=>X"0000045700000458000004590000045a", 2106=>X"00000452000004530000045400000456", 2107=>X"0000044d0000044f0000045000000451", 2108=>X"000004490000044a0000044b0000044c", 2109=>X"00000444000004450000044700000448", 
2110=>X"00000440000004410000044200000443", 2111=>X"0000043b0000043c0000043d0000043f", 2112=>X"0000043700000438000004390000043a", 2113=>X"00000432000004330000043500000436", 2114=>X"0000042e0000042f0000043000000431", 
2115=>X"0000042a0000042b0000042c0000042d", 2116=>X"00000425000004260000042700000429", 2117=>X"00000421000004220000042300000424", 2118=>X"0000041d0000041e0000041f00000420", 2119=>X"000004190000041a0000041b0000041c", 
2120=>X"00000414000004150000041600000418", 2121=>X"00000410000004110000041200000413", 2122=>X"0000040c0000040d0000040e0000040f", 2123=>X"00000408000004090000040a0000040b", 2124=>X"00000404000004050000040600000407", 
2125=>X"00000400000004010000040200000403", 2126=>X"000003fc000003fd000003fe000003ff", 2127=>X"000003f8000003f9000003fa000003fb", 2128=>X"000003f4000003f5000003f6000003f7", 2129=>X"000003f0000003f1000003f2000003f3", 
2130=>X"000003ec000003ed000003ee000003ef", 2131=>X"000003e9000003ea000003ea000003eb", 2132=>X"000003e5000003e6000003e7000003e8", 2133=>X"000003e1000003e2000003e3000003e4", 2134=>X"000003dd000003de000003df000003e0", 
2135=>X"000003da000003da000003db000003dc", 2136=>X"000003d6000003d7000003d8000003d9", 2137=>X"000003d2000003d3000003d4000003d5", 2138=>X"000003cf000003cf000003d0000003d1", 2139=>X"000003cb000003cc000003cd000003ce", 
2140=>X"000003c7000003c8000003c9000003ca", 2141=>X"000003c4000003c5000003c6000003c6", 2142=>X"000003c0000003c1000003c2000003c3", 2143=>X"000003bd000003be000003be000003bf", 2144=>X"000003b9000003ba000003bb000003bc", 
2145=>X"000003b6000003b7000003b8000003b8", 2146=>X"000003b2000003b3000003b4000003b5", 2147=>X"000003af000003b0000003b1000003b2", 2148=>X"000003ac000003ac000003ad000003ae", 2149=>X"000003a8000003a9000003aa000003ab", 
2150=>X"000003a5000003a6000003a7000003a7", 2151=>X"000003a2000003a2000003a3000003a4", 2152=>X"0000039e0000039f000003a0000003a1", 2153=>X"0000039b0000039c0000039d0000039d", 2154=>X"0000039800000399000003990000039a", 
2155=>X"00000395000003950000039600000397", 2156=>X"00000391000003920000039300000394", 2157=>X"0000038e0000038f0000039000000391", 2158=>X"0000038b0000038c0000038d0000038d", 2159=>X"00000388000003890000038a0000038a", 
2160=>X"00000385000003860000038600000387", 2161=>X"00000382000003830000038300000384", 2162=>X"0000037f0000037f0000038000000381", 2163=>X"0000037c0000037c0000037d0000037e", 2164=>X"00000379000003790000037a0000037b", 
2165=>X"00000376000003760000037700000378", 2166=>X"00000373000003730000037400000375", 2167=>X"00000370000003700000037100000372", 2168=>X"0000036d0000036d0000036e0000036f", 2169=>X"0000036a0000036b0000036b0000036c", 
2170=>X"00000367000003680000036800000369", 2171=>X"00000364000003650000036500000366", 2172=>X"00000361000003620000036300000363", 2173=>X"0000035e0000035f0000036000000360", 2174=>X"0000035b0000035c0000035d0000035e", 
2175=>X"00000359000003590000035a0000035b", 2176=>X"00000356000003570000035700000358", 2177=>X"00000353000003540000035500000355", 2178=>X"00000350000003510000035200000352", 2179=>X"0000034e0000034e0000034f00000350", 
2180=>X"0000034b0000034c0000034c0000034d", 2181=>X"00000348000003490000034a0000034a", 2182=>X"00000346000003460000034700000348", 2183=>X"00000343000003440000034400000345", 2184=>X"00000340000003410000034200000342", 
2185=>X"0000033e0000033e0000033f00000340", 2186=>X"0000033b0000033c0000033c0000033d", 2187=>X"00000338000003390000033a0000033a", 2188=>X"00000336000003360000033700000338", 2189=>X"00000333000003340000033400000335", 
2190=>X"00000331000003310000033200000333", 2191=>X"0000032e0000032f0000032f00000330", 2192=>X"0000032c0000032c0000032d0000032d", 2193=>X"000003290000032a0000032a0000032b", 2194=>X"00000327000003270000032800000328", 
2195=>X"00000324000003250000032500000326", 2196=>X"00000322000003220000032300000324", 2197=>X"0000031f000003200000032000000321", 2198=>X"0000031d0000031d0000031e0000031f", 2199=>X"0000031a0000031b0000031c0000031c", 
2200=>X"0000031800000319000003190000031a", 2201=>X"00000316000003160000031700000317", 2202=>X"00000313000003140000031400000315", 2203=>X"00000311000003110000031200000313", 2204=>X"0000030f0000030f0000031000000310", 
2205=>X"0000030c0000030d0000030d0000030e", 2206=>X"0000030a0000030a0000030b0000030c", 2207=>X"00000308000003080000030900000309", 2208=>X"00000305000003060000030600000307", 2209=>X"00000303000003040000030400000305", 
2210=>X"00000301000003010000030200000302", 2211=>X"000002ff000002ff0000030000000300", 2212=>X"000002fc000002fd000002fd000002fe", 2213=>X"000002fa000002fb000002fb000002fc", 2214=>X"000002f8000002f8000002f9000002f9", 
2215=>X"000002f6000002f6000002f7000002f7", 2216=>X"000002f3000002f4000002f5000002f5", 2217=>X"000002f1000002f2000002f2000002f3", 2218=>X"000002ef000002f0000002f0000002f1", 2219=>X"000002ed000002ee000002ee000002ef", 
2220=>X"000002eb000002eb000002ec000002ec", 2221=>X"000002e9000002e9000002ea000002ea", 2222=>X"000002e7000002e7000002e8000002e8", 2223=>X"000002e5000002e5000002e6000002e6", 2224=>X"000002e2000002e3000002e3000002e4", 
2225=>X"000002e0000002e1000002e1000002e2", 2226=>X"000002de000002df000002df000002e0", 2227=>X"000002dc000002dd000002dd000002de", 2228=>X"000002da000002db000002db000002dc", 2229=>X"000002d8000002d9000002d9000002da", 
2230=>X"000002d6000002d7000002d7000002d8", 2231=>X"000002d4000002d5000002d5000002d6", 2232=>X"000002d2000002d3000002d3000002d4", 2233=>X"000002d0000002d1000002d1000002d2", 2234=>X"000002ce000002cf000002cf000002d0", 
2235=>X"000002cc000002cd000002cd000002ce", 2236=>X"000002ca000002cb000002cb000002cc", 2237=>X"000002c8000002c9000002c9000002ca", 2238=>X"000002c6000002c7000002c7000002c8", 2239=>X"000002c4000002c5000002c5000002c6", 
2240=>X"000002c3000002c3000002c4000002c4", 2241=>X"000002c1000002c1000002c2000002c2", 2242=>X"000002bf000002bf000002c0000002c0", 2243=>X"000002bd000002bd000002be000002be", 2244=>X"000002bb000002bc000002bc000002bc", 
2245=>X"000002b9000002ba000002ba000002bb", 2246=>X"000002b7000002b8000002b8000002b9", 2247=>X"000002b6000002b6000002b6000002b7", 2248=>X"000002b4000002b4000002b5000002b5", 2249=>X"000002b2000002b2000002b3000002b3", 
2250=>X"000002b0000002b0000002b1000002b1", 2251=>X"000002ae000002af000002af000002b0", 2252=>X"000002ac000002ad000002ad000002ae", 2253=>X"000002ab000002ab000002ac000002ac", 2254=>X"000002a9000002a9000002aa000002aa", 
2255=>X"000002a7000002a8000002a8000002a8", 2256=>X"000002a5000002a6000002a6000002a7", 2257=>X"000002a4000002a4000002a5000002a5", 2258=>X"000002a2000002a2000002a3000002a3", 2259=>X"000002a0000002a1000002a1000002a1", 
2260=>X"0000029e0000029f0000029f000002a0", 2261=>X"0000029d0000029d0000029e0000029e", 2262=>X"0000029b0000029b0000029c0000029c", 2263=>X"000002990000029a0000029a0000029b", 2264=>X"00000298000002980000029800000299", 
2265=>X"00000296000002960000029700000297", 2266=>X"00000294000002950000029500000296", 2267=>X"00000293000002930000029300000294", 2268=>X"00000291000002910000029200000292", 2269=>X"0000028f000002900000029000000291", 
2270=>X"0000028e0000028e0000028f0000028f", 2271=>X"0000028c0000028d0000028d0000028d", 2272=>X"0000028a0000028b0000028b0000028c", 2273=>X"00000289000002890000028a0000028a", 2274=>X"00000287000002880000028800000288", 
2275=>X"00000286000002860000028600000287", 2276=>X"00000284000002840000028500000285", 2277=>X"00000283000002830000028300000284", 2278=>X"00000281000002810000028200000282", 2279=>X"0000027f000002800000028000000281", 
2280=>X"0000027e0000027e0000027f0000027f", 2281=>X"0000027c0000027d0000027d0000027d", 2282=>X"0000027b0000027b0000027c0000027c", 2283=>X"000002790000027a0000027a0000027a", 2284=>X"00000278000002780000027800000279", 
2285=>X"00000276000002770000027700000277", 2286=>X"00000275000002750000027500000276", 2287=>X"00000273000002740000027400000274", 2288=>X"00000272000002720000027200000273", 2289=>X"00000270000002710000027100000271", 
2290=>X"0000026f0000026f0000026f00000270", 2291=>X"0000026d0000026e0000026e0000026e", 2292=>X"0000026c0000026c0000026c0000026d", 2293=>X"0000026a0000026b0000026b0000026b", 2294=>X"00000269000002690000026a0000026a", 
2295=>X"00000267000002680000026800000268", 2296=>X"00000266000002660000026700000267", 2297=>X"00000264000002650000026500000266", 2298=>X"00000263000002630000026400000264", 2299=>X"00000262000002620000026200000263", 
2300=>X"00000260000002610000026100000261", 2301=>X"0000025f0000025f0000026000000260", 2302=>X"0000025d0000025e0000025e0000025e", 2303=>X"0000025c0000025c0000025d0000025d", 2304=>X"0000025b0000025b0000025b0000025c", 
2305=>X"000002590000025a0000025a0000025a", 2306=>X"00000258000002580000025900000259", 2307=>X"00000257000002570000025700000258", 2308=>X"00000255000002550000025600000256", 2309=>X"00000254000002540000025400000255", 
2310=>X"00000252000002530000025300000253", 2311=>X"00000251000002510000025200000252", 2312=>X"00000250000002500000025000000251", 2313=>X"0000024e0000024f0000024f0000024f", 2314=>X"0000024d0000024d0000024e0000024e", 
2315=>X"0000024c0000024c0000024c0000024d", 2316=>X"0000024a0000024b0000024b0000024b", 2317=>X"00000249000002490000024a0000024a", 2318=>X"00000248000002480000024800000249", 2319=>X"00000247000002470000024700000248", 
2320=>X"00000245000002460000024600000246", 2321=>X"00000244000002440000024500000245", 2322=>X"00000243000002430000024300000244", 2323=>X"00000241000002420000024200000242", 2324=>X"00000240000002400000024100000241", 
2325=>X"0000023f0000023f0000024000000240", 2326=>X"0000023e0000023e0000023e0000023f", 2327=>X"0000023c0000023d0000023d0000023d", 2328=>X"0000023b0000023b0000023c0000023c", 2329=>X"0000023a0000023a0000023a0000023b", 
2330=>X"0000023900000239000002390000023a", 2331=>X"00000237000002380000023800000238", 2332=>X"00000236000002360000023700000237", 2333=>X"00000235000002350000023600000236", 2334=>X"00000234000002340000023400000235", 
2335=>X"00000233000002330000023300000233", 2336=>X"00000231000002320000023200000232", 2337=>X"00000230000002300000023100000231", 2338=>X"0000022f0000022f0000023000000230", 2339=>X"0000022e0000022e0000022e0000022f", 
2340=>X"0000022d0000022d0000022d0000022d", 2341=>X"0000022b0000022c0000022c0000022c", 2342=>X"0000022a0000022b0000022b0000022b", 2343=>X"00000229000002290000022a0000022a", 2344=>X"00000228000002280000022800000229", 
2345=>X"00000227000002270000022700000228", 2346=>X"00000226000002260000022600000226", 2347=>X"00000224000002250000022500000225", 2348=>X"00000223000002240000022400000224", 2349=>X"00000222000002220000022300000223", 
2350=>X"00000221000002210000022200000222", 2351=>X"00000220000002200000022000000221", 2352=>X"0000021f0000021f0000021f00000220", 2353=>X"0000021e0000021e0000021e0000021e", 2354=>X"0000021d0000021d0000021d0000021d", 
2355=>X"0000021b0000021c0000021c0000021c", 2356=>X"0000021a0000021b0000021b0000021b", 2357=>X"00000219000002190000021a0000021a", 2358=>X"00000218000002180000021900000219", 2359=>X"00000217000002170000021800000218", 
2360=>X"00000216000002160000021600000217", 2361=>X"00000215000002150000021500000216", 2362=>X"00000214000002140000021400000215", 2363=>X"00000213000002130000021300000213", 2364=>X"00000212000002120000021200000212", 
2365=>X"00000211000002110000021100000211", 2366=>X"0000020f000002100000021000000210", 2367=>X"0000020e0000020f0000020f0000020f", 2368=>X"0000020d0000020e0000020e0000020e", 2369=>X"0000020c0000020d0000020d0000020d", 
2370=>X"0000020b0000020c0000020c0000020c", 2371=>X"0000020a0000020a0000020b0000020b", 2372=>X"00000209000002090000020a0000020a", 2373=>X"00000208000002080000020900000209", 2374=>X"00000207000002070000020800000208", 
2375=>X"00000206000002060000020700000207", 2376=>X"00000205000002050000020600000206", 2377=>X"00000204000002040000020500000205", 2378=>X"00000203000002030000020400000204", 2379=>X"00000202000002020000020300000203", 
2380=>X"00000201000002010000020200000202", 2381=>X"00000200000002000000020100000201", 2382=>X"000001ff000001ff0000020000000200", 2383=>X"000001fe000001fe000001ff000001ff", 2384=>X"000001fd000001fd000001fe000001fe", 
2385=>X"000001fc000001fc000001fd000001fd", 2386=>X"000001fb000001fb000001fc000001fc", 2387=>X"000001fa000001fa000001fb000001fb", 2388=>X"000001f9000001f9000001fa000001fa", 2389=>X"000001f8000001f8000001f9000001f9", 
2390=>X"000001f7000001f7000001f8000001f8", 2391=>X"000001f6000001f6000001f7000001f7", 2392=>X"000001f5000001f5000001f6000001f6", 2393=>X"000001f4000001f5000001f5000001f5", 2394=>X"000001f3000001f4000001f4000001f4", 
2395=>X"000001f2000001f3000001f3000001f3", 2396=>X"000001f1000001f2000001f2000001f2", 2397=>X"000001f0000001f1000001f1000001f1", 2398=>X"000001f0000001f0000001f0000001f0", 2399=>X"000001ef000001ef000001ef000001ef", 
2400=>X"000001ee000001ee000001ee000001ee", 2401=>X"000001ed000001ed000001ed000001ed", 2402=>X"000001ec000001ec000001ec000001ed", 2403=>X"000001eb000001eb000001eb000001ec", 2404=>X"000001ea000001ea000001ea000001eb", 
2405=>X"000001e9000001e9000001ea000001ea", 2406=>X"000001e8000001e8000001e9000001e9", 2407=>X"000001e7000001e7000001e8000001e8", 2408=>X"000001e6000001e7000001e7000001e7", 2409=>X"000001e5000001e6000001e6000001e6", 
2410=>X"000001e5000001e5000001e5000001e5", 2411=>X"000001e4000001e4000001e4000001e4", 2412=>X"000001e3000001e3000001e3000001e3", 2413=>X"000001e2000001e2000001e2000001e3", 2414=>X"000001e1000001e1000001e1000001e2", 
2415=>X"000001e0000001e0000001e1000001e1", 2416=>X"000001df000001df000001e0000001e0", 2417=>X"000001de000001df000001df000001df", 2418=>X"000001dd000001de000001de000001de", 2419=>X"000001dd000001dd000001dd000001dd", 
2420=>X"000001dc000001dc000001dc000001dc", 2421=>X"000001db000001db000001db000001dc", 2422=>X"000001da000001da000001da000001db", 2423=>X"000001d9000001d9000001da000001da", 2424=>X"000001d8000001d9000001d9000001d9", 
2425=>X"000001d7000001d8000001d8000001d8", 2426=>X"000001d7000001d7000001d7000001d7", 2427=>X"000001d6000001d6000001d6000001d6", 2428=>X"000001d5000001d5000001d5000001d6", 2429=>X"000001d4000001d4000001d5000001d5", 
2430=>X"000001d3000001d3000001d4000001d4", 2431=>X"000001d2000001d3000001d3000001d3", 2432=>X"000001d2000001d2000001d2000001d2", 2433=>X"000001d1000001d1000001d1000001d1", 2434=>X"000001d0000001d0000001d0000001d1", 
2435=>X"000001cf000001cf000001d0000001d0", 2436=>X"000001ce000001cf000001cf000001cf", 2437=>X"000001ce000001ce000001ce000001ce", 2438=>X"000001cd000001cd000001cd000001cd", 2439=>X"000001cc000001cc000001cc000001cd", 
2440=>X"000001cb000001cb000001cb000001cc", 2441=>X"000001ca000001ca000001cb000001cb", 2442=>X"000001c9000001ca000001ca000001ca", 2443=>X"000001c9000001c9000001c9000001c9", 2444=>X"000001c8000001c8000001c8000001c8", 
2445=>X"000001c7000001c7000001c8000001c8", 2446=>X"000001c6000001c7000001c7000001c7", 2447=>X"000001c6000001c6000001c6000001c6", 2448=>X"000001c5000001c5000001c5000001c5", 2449=>X"000001c4000001c4000001c4000001c5", 
2450=>X"000001c3000001c3000001c4000001c4", 2451=>X"000001c2000001c3000001c3000001c3", 2452=>X"000001c2000001c2000001c2000001c2", 2453=>X"000001c1000001c1000001c1000001c1", 2454=>X"000001c0000001c0000001c0000001c1", 
2455=>X"000001bf000001c0000001c0000001c0", 2456=>X"000001bf000001bf000001bf000001bf", 2457=>X"000001be000001be000001be000001be", 2458=>X"000001bd000001bd000001bd000001be", 2459=>X"000001bc000001bd000001bd000001bd", 
2460=>X"000001bc000001bc000001bc000001bc", 2461=>X"000001bb000001bb000001bb000001bb", 2462=>X"000001ba000001ba000001ba000001bb", 2463=>X"000001b9000001ba000001ba000001ba", 2464=>X"000001b9000001b9000001b9000001b9", 
2465=>X"000001b8000001b8000001b8000001b8", 2466=>X"000001b7000001b7000001b7000001b8", 2467=>X"000001b6000001b7000001b7000001b7", 2468=>X"000001b6000001b6000001b6000001b6", 2469=>X"000001b5000001b5000001b5000001b5", 
2470=>X"000001b4000001b4000001b5000001b5", 2471=>X"000001b3000001b4000001b4000001b4", 2472=>X"000001b3000001b3000001b3000001b3", 2473=>X"000001b2000001b2000001b2000001b3", 2474=>X"000001b1000001b1000001b2000001b2", 
2475=>X"000001b1000001b1000001b1000001b1", 2476=>X"000001b0000001b0000001b0000001b0", 2477=>X"000001af000001af000001b0000001b0", 2478=>X"000001ae000001af000001af000001af", 2479=>X"000001ae000001ae000001ae000001ae", 
2480=>X"000001ad000001ad000001ad000001ae", 2481=>X"000001ac000001ad000001ad000001ad", 2482=>X"000001ac000001ac000001ac000001ac", 2483=>X"000001ab000001ab000001ab000001ab", 2484=>X"000001aa000001aa000001ab000001ab", 
2485=>X"000001aa000001aa000001aa000001aa", 2486=>X"000001a9000001a9000001a9000001a9", 2487=>X"000001a8000001a8000001a9000001a9", 2488=>X"000001a7000001a8000001a8000001a8", 2489=>X"000001a7000001a7000001a7000001a7", 
2490=>X"000001a6000001a6000001a6000001a7", 2491=>X"000001a5000001a6000001a6000001a6", 2492=>X"000001a5000001a5000001a5000001a5", 2493=>X"000001a4000001a4000001a4000001a5", 2494=>X"000001a3000001a4000001a4000001a4", 
2495=>X"000001a3000001a3000001a3000001a3", 2496=>X"000001a2000001a2000001a2000001a3", 2497=>X"000001a1000001a2000001a2000001a2", 2498=>X"000001a1000001a1000001a1000001a1", 2499=>X"000001a0000001a0000001a0000001a1", 
2500=>X"0000019f000001a0000001a0000001a0", 2501=>X"0000019f0000019f0000019f0000019f", 2502=>X"0000019e0000019e0000019e0000019f", 2503=>X"0000019d0000019e0000019e0000019e", 2504=>X"0000019d0000019d0000019d0000019d", 
2505=>X"0000019c0000019c0000019d0000019d", 2506=>X"0000019c0000019c0000019c0000019c", 2507=>X"0000019b0000019b0000019b0000019b", 2508=>X"0000019a0000019a0000019b0000019b", 2509=>X"0000019a0000019a0000019a0000019a", 
2510=>X"00000199000001990000019900000199", 2511=>X"00000198000001980000019900000199", 2512=>X"00000198000001980000019800000198", 2513=>X"00000197000001970000019700000198", 2514=>X"00000196000001970000019700000197", 
2515=>X"00000196000001960000019600000196", 2516=>X"00000195000001950000019500000196", 2517=>X"00000195000001950000019500000195", 2518=>X"00000194000001940000019400000194", 2519=>X"00000193000001930000019400000194", 
2520=>X"00000193000001930000019300000193", 2521=>X"00000192000001920000019200000193", 2522=>X"00000191000001920000019200000192", 2523=>X"00000191000001910000019100000191", 2524=>X"00000190000001900000019100000191", 
2525=>X"00000190000001900000019000000190", 2526=>X"0000018f0000018f0000018f0000018f", 2527=>X"0000018e0000018f0000018f0000018f", 2528=>X"0000018e0000018e0000018e0000018e", 2529=>X"0000018d0000018d0000018d0000018e", 
2530=>X"0000018d0000018d0000018d0000018d", 2531=>X"0000018c0000018c0000018c0000018c", 2532=>X"0000018b0000018c0000018c0000018c", 2533=>X"0000018b0000018b0000018b0000018b", 2534=>X"0000018a0000018a0000018a0000018b", 
2535=>X"0000018a0000018a0000018a0000018a", 2536=>X"00000189000001890000018900000189", 2537=>X"00000188000001890000018900000189", 2538=>X"00000188000001880000018800000188", 2539=>X"00000187000001870000018800000188", 
2540=>X"00000187000001870000018700000187", 2541=>X"00000186000001860000018600000187", 2542=>X"00000186000001860000018600000186", 2543=>X"00000185000001850000018500000185", 2544=>X"00000184000001850000018500000185", 
2545=>X"00000184000001840000018400000184", 2546=>X"00000183000001830000018400000184", 2547=>X"00000183000001830000018300000183", 2548=>X"00000182000001820000018200000183", 2549=>X"00000182000001820000018200000182", 
2550=>X"00000181000001810000018100000181", 2551=>X"00000180000001810000018100000181", 2552=>X"00000180000001800000018000000180", 2553=>X"0000017f0000017f0000018000000180", 2554=>X"0000017f0000017f0000017f0000017f", 
2555=>X"0000017e0000017e0000017e0000017f", 2556=>X"0000017e0000017e0000017e0000017e", 2557=>X"0000017d0000017d0000017d0000017d", 2558=>X"0000017c0000017d0000017d0000017d", 2559=>X"0000017c0000017c0000017c0000017c", 
2560=>X"0000017b0000017c0000017c0000017c", 2561=>X"0000017b0000017b0000017b0000017b", 2562=>X"0000017a0000017a0000017b0000017b", 2563=>X"0000017a0000017a0000017a0000017a", 2564=>X"0000017900000179000001790000017a", 
2565=>X"00000179000001790000017900000179", 2566=>X"00000178000001780000017800000179", 2567=>X"00000178000001780000017800000178", 2568=>X"00000177000001770000017700000177", 2569=>X"00000176000001770000017700000177", 
2570=>X"00000176000001760000017600000176", 2571=>X"00000175000001760000017600000176", 2572=>X"00000175000001750000017500000175", 2573=>X"00000174000001740000017500000175", 2574=>X"00000174000001740000017400000174", 
2575=>X"00000173000001730000017400000174", 2576=>X"00000173000001730000017300000173", 2577=>X"00000172000001720000017300000173", 2578=>X"00000172000001720000017200000172", 2579=>X"00000171000001710000017100000172", 
2580=>X"00000171000001710000017100000171", 2581=>X"00000170000001700000017000000171", 2582=>X"00000170000001700000017000000170", 2583=>X"0000016f0000016f0000016f00000170", 2584=>X"0000016f0000016f0000016f0000016f", 
2585=>X"0000016e0000016e0000016e0000016f", 2586=>X"0000016e0000016e0000016e0000016e", 2587=>X"0000016d0000016d0000016d0000016d", 2588=>X"0000016d0000016d0000016d0000016d", 2589=>X"0000016c0000016c0000016c0000016c", 
2590=>X"0000016c0000016c0000016c0000016c", 2591=>X"0000016b0000016b0000016b0000016b", 2592=>X"0000016b0000016b0000016b0000016b", 2593=>X"0000016a0000016a0000016a0000016a", 2594=>X"0000016a0000016a0000016a0000016a", 
2595=>X"00000169000001690000016900000169", 2596=>X"00000169000001690000016900000169", 2597=>X"00000168000001680000016800000168", 2598=>X"00000168000001680000016800000168", 2599=>X"00000167000001670000016700000167", 
2600=>X"00000167000001670000016700000167", 2601=>X"00000166000001660000016600000166", 2602=>X"00000166000001660000016600000166", 2603=>X"00000165000001650000016500000166", 2604=>X"00000165000001650000016500000165", 
2605=>X"00000164000001640000016400000165", 2606=>X"00000164000001640000016400000164", 2607=>X"00000163000001630000016300000164", 2608=>X"00000163000001630000016300000163", 2609=>X"00000162000001620000016200000163", 
2610=>X"00000162000001620000016200000162", 2611=>X"00000161000001610000016200000162", 2612=>X"00000161000001610000016100000161", 2613=>X"00000160000001600000016100000161", 2614=>X"00000160000001600000016000000160", 
2615=>X"0000015f000001600000016000000160", 2616=>X"0000015f0000015f0000015f0000015f", 2617=>X"0000015e0000015f0000015f0000015f", 2618=>X"0000015e0000015e0000015e0000015e", 2619=>X"0000015e0000015e0000015e0000015e", 
2620=>X"0000015d0000015d0000015d0000015d", 2621=>X"0000015d0000015d0000015d0000015d", 2622=>X"0000015c0000015c0000015c0000015c", 2623=>X"0000015c0000015c0000015c0000015c", 2624=>X"0000015b0000015b0000015b0000015c", 
2625=>X"0000015b0000015b0000015b0000015b", 2626=>X"0000015a0000015a0000015b0000015b", 2627=>X"0000015a0000015a0000015a0000015a", 2628=>X"00000159000001590000015a0000015a", 2629=>X"00000159000001590000015900000159", 
2630=>X"00000158000001590000015900000159", 2631=>X"00000158000001580000015800000158", 2632=>X"00000158000001580000015800000158", 2633=>X"00000157000001570000015700000157", 2634=>X"00000157000001570000015700000157", 
2635=>X"00000156000001560000015600000157", 2636=>X"00000156000001560000015600000156", 2637=>X"00000155000001550000015600000156", 2638=>X"00000155000001550000015500000155", 2639=>X"00000154000001550000015500000155", 
2640=>X"00000154000001540000015400000154", 2641=>X"00000154000001540000015400000154", 2642=>X"00000153000001530000015300000153", 2643=>X"00000153000001530000015300000153", 2644=>X"00000152000001520000015200000153", 
2645=>X"00000152000001520000015200000152", 2646=>X"00000151000001510000015200000152", 2647=>X"00000151000001510000015100000151", 2648=>X"00000151000001510000015100000151", 2649=>X"00000150000001500000015000000150", 
2650=>X"00000150000001500000015000000150", 2651=>X"0000014f0000014f0000014f00000150", 2652=>X"0000014f0000014f0000014f0000014f", 2653=>X"0000014e0000014e0000014f0000014f", 2654=>X"0000014e0000014e0000014e0000014e", 
2655=>X"0000014e0000014e0000014e0000014e", 2656=>X"0000014d0000014d0000014d0000014d", 2657=>X"0000014d0000014d0000014d0000014d", 2658=>X"0000014c0000014c0000014c0000014d", 2659=>X"0000014c0000014c0000014c0000014c", 
2660=>X"0000014b0000014c0000014c0000014c", 2661=>X"0000014b0000014b0000014b0000014b", 2662=>X"0000014b0000014b0000014b0000014b", 2663=>X"0000014a0000014a0000014a0000014a", 2664=>X"0000014a0000014a0000014a0000014a", 
2665=>X"00000149000001490000014a0000014a", 2666=>X"00000149000001490000014900000149", 2667=>X"00000149000001490000014900000149", 2668=>X"00000148000001480000014800000148", 2669=>X"00000148000001480000014800000148", 
2670=>X"00000147000001470000014700000148", 2671=>X"00000147000001470000014700000147", 2672=>X"00000146000001470000014700000147", 2673=>X"00000146000001460000014600000146", 2674=>X"00000146000001460000014600000146", 
2675=>X"00000145000001450000014500000146", 2676=>X"00000145000001450000014500000145", 2677=>X"00000144000001450000014500000145", 2678=>X"00000144000001440000014400000144", 2679=>X"00000144000001440000014400000144", 
2680=>X"00000143000001430000014300000144", 2681=>X"00000143000001430000014300000143", 2682=>X"00000142000001430000014300000143", 2683=>X"00000142000001420000014200000142", 2684=>X"00000142000001420000014200000142", 
2685=>X"00000141000001410000014100000142", 2686=>X"00000141000001410000014100000141", 2687=>X"00000140000001410000014100000141", 2688=>X"00000140000001400000014000000140", 2689=>X"00000140000001400000014000000140", 
2690=>X"0000013f0000013f0000013f00000140", 2691=>X"0000013f0000013f0000013f0000013f", 2692=>X"0000013f0000013f0000013f0000013f", 2693=>X"0000013e0000013e0000013e0000013e", 2694=>X"0000013e0000013e0000013e0000013e", 
2695=>X"0000013d0000013d0000013e0000013e", 2696=>X"0000013d0000013d0000013d0000013d", 2697=>X"0000013d0000013d0000013d0000013d", 2698=>X"0000013c0000013c0000013c0000013d", 2699=>X"0000013c0000013c0000013c0000013c", 
2700=>X"0000013b0000013c0000013c0000013c", 2701=>X"0000013b0000013b0000013b0000013b", 2702=>X"0000013b0000013b0000013b0000013b", 2703=>X"0000013a0000013a0000013b0000013b", 2704=>X"0000013a0000013a0000013a0000013a", 
2705=>X"0000013a0000013a0000013a0000013a", 2706=>X"00000139000001390000013900000139", 2707=>X"00000139000001390000013900000139", 2708=>X"00000138000001390000013900000139", 2709=>X"00000138000001380000013800000138", 
2710=>X"00000138000001380000013800000138", 2711=>X"00000137000001370000013800000138", 2712=>X"00000137000001370000013700000137", 2713=>X"00000137000001370000013700000137", 2714=>X"00000136000001360000013600000137", 
2715=>X"00000136000001360000013600000136", 2716=>X"00000135000001360000013600000136", 2717=>X"00000135000001350000013500000135", 2718=>X"00000135000001350000013500000135", 2719=>X"00000134000001340000013500000135", 
2720=>X"00000134000001340000013400000134", 2721=>X"00000134000001340000013400000134", 2722=>X"00000133000001330000013400000134", 2723=>X"00000133000001330000013300000133", 2724=>X"00000133000001330000013300000133", 
2725=>X"00000132000001320000013200000133", 2726=>X"00000132000001320000013200000132", 2727=>X"00000132000001320000013200000132", 2728=>X"00000131000001310000013100000131", 2729=>X"00000131000001310000013100000131", 
2730=>X"00000130000001310000013100000131", 2731=>X"00000130000001300000013000000130", 2732=>X"00000130000001300000013000000130", 2733=>X"0000012f0000012f0000013000000130", 2734=>X"0000012f0000012f0000012f0000012f", 
2735=>X"0000012f0000012f0000012f0000012f", 2736=>X"0000012e0000012e0000012f0000012f", 2737=>X"0000012e0000012e0000012e0000012e", 2738=>X"0000012e0000012e0000012e0000012e", 2739=>X"0000012d0000012d0000012d0000012e", 
2740=>X"0000012d0000012d0000012d0000012d", 2741=>X"0000012d0000012d0000012d0000012d", 2742=>X"0000012c0000012c0000012c0000012d", 2743=>X"0000012c0000012c0000012c0000012c", 2744=>X"0000012c0000012c0000012c0000012c", 
2745=>X"0000012b0000012b0000012b0000012c", 2746=>X"0000012b0000012b0000012b0000012b", 2747=>X"0000012b0000012b0000012b0000012b", 2748=>X"0000012a0000012a0000012a0000012a", 2749=>X"0000012a0000012a0000012a0000012a", 
2750=>X"0000012a0000012a0000012a0000012a", 2751=>X"00000129000001290000012900000129", 2752=>X"00000129000001290000012900000129", 2753=>X"00000129000001290000012900000129", 2754=>X"00000128000001280000012800000128", 
2755=>X"00000128000001280000012800000128", 2756=>X"00000128000001280000012800000128", 2757=>X"00000127000001270000012700000127", 2758=>X"00000127000001270000012700000127", 2759=>X"00000127000001270000012700000127", 
2760=>X"00000126000001260000012600000126", 2761=>X"00000126000001260000012600000126", 2762=>X"00000126000001260000012600000126", 2763=>X"00000125000001250000012500000125", 2764=>X"00000125000001250000012500000125", 
2765=>X"00000125000001250000012500000125", 2766=>X"00000124000001240000012400000124", 2767=>X"00000124000001240000012400000124", 2768=>X"00000124000001240000012400000124", 2769=>X"00000123000001230000012300000124", 
2770=>X"00000123000001230000012300000123", 2771=>X"00000123000001230000012300000123", 2772=>X"00000122000001220000012200000123", 2773=>X"00000122000001220000012200000122", 2774=>X"00000122000001220000012200000122", 
2775=>X"00000121000001210000012200000122", 2776=>X"00000121000001210000012100000121", 2777=>X"00000121000001210000012100000121", 2778=>X"00000120000001200000012100000121", 2779=>X"00000120000001200000012000000120", 
2780=>X"00000120000001200000012000000120", 2781=>X"0000011f000001200000012000000120", 2782=>X"0000011f0000011f0000011f0000011f", 2783=>X"0000011f0000011f0000011f0000011f", 2784=>X"0000011e0000011f0000011f0000011f", 
2785=>X"0000011e0000011e0000011e0000011e", 2786=>X"0000011e0000011e0000011e0000011e", 2787=>X"0000011e0000011e0000011e0000011e", 2788=>X"0000011d0000011d0000011d0000011d", 2789=>X"0000011d0000011d0000011d0000011d", 
2790=>X"0000011d0000011d0000011d0000011d", 2791=>X"0000011c0000011c0000011c0000011d", 2792=>X"0000011c0000011c0000011c0000011c", 2793=>X"0000011c0000011c0000011c0000011c", 2794=>X"0000011b0000011b0000011c0000011c", 
2795=>X"0000011b0000011b0000011b0000011b", 2796=>X"0000011b0000011b0000011b0000011b", 2797=>X"0000011a0000011b0000011b0000011b", 2798=>X"0000011a0000011a0000011a0000011a", 2799=>X"0000011a0000011a0000011a0000011a", 
2800=>X"0000011a0000011a0000011a0000011a", 2801=>X"00000119000001190000011900000119", 2802=>X"00000119000001190000011900000119", 2803=>X"00000119000001190000011900000119", 2804=>X"00000118000001180000011900000119", 
2805=>X"00000118000001180000011800000118", 2806=>X"00000118000001180000011800000118", 2807=>X"00000117000001180000011800000118", 2808=>X"00000117000001170000011700000117", 2809=>X"00000117000001170000011700000117", 
2810=>X"00000117000001170000011700000117", 2811=>X"00000116000001160000011600000117", 2812=>X"00000116000001160000011600000116", 2813=>X"00000116000001160000011600000116", 2814=>X"00000115000001150000011600000116", 
2815=>X"00000115000001150000011500000115", 2816=>X"00000115000001150000011500000115", 2817=>X"00000115000001150000011500000115", 2818=>X"00000114000001140000011400000114", 2819=>X"00000114000001140000011400000114", 
2820=>X"00000114000001140000011400000114", 2821=>X"00000113000001130000011400000114", 2822=>X"00000113000001130000011300000113", 2823=>X"00000113000001130000011300000113", 2824=>X"00000112000001130000011300000113", 
2825=>X"00000112000001120000011200000112", 2826=>X"00000112000001120000011200000112", 2827=>X"00000112000001120000011200000112", 2828=>X"00000111000001110000011100000112", 2829=>X"00000111000001110000011100000111", 
2830=>X"00000111000001110000011100000111", 2831=>X"00000110000001110000011100000111", 2832=>X"00000110000001100000011000000110", 2833=>X"00000110000001100000011000000110", 2834=>X"00000110000001100000011000000110", 
2835=>X"0000010f0000010f0000011000000110", 2836=>X"0000010f0000010f0000010f0000010f", 2837=>X"0000010f0000010f0000010f0000010f", 2838=>X"0000010f0000010f0000010f0000010f", 2839=>X"0000010e0000010e0000010e0000010e", 
2840=>X"0000010e0000010e0000010e0000010e", 2841=>X"0000010e0000010e0000010e0000010e", 2842=>X"0000010d0000010d0000010e0000010e", 2843=>X"0000010d0000010d0000010d0000010d", 2844=>X"0000010d0000010d0000010d0000010d", 
2845=>X"0000010d0000010d0000010d0000010d", 2846=>X"0000010c0000010c0000010c0000010d", 2847=>X"0000010c0000010c0000010c0000010c", 2848=>X"0000010c0000010c0000010c0000010c", 2849=>X"0000010b0000010c0000010c0000010c", 
2850=>X"0000010b0000010b0000010b0000010b", 2851=>X"0000010b0000010b0000010b0000010b", 2852=>X"0000010b0000010b0000010b0000010b", 2853=>X"0000010a0000010a0000010b0000010b", 2854=>X"0000010a0000010a0000010a0000010a", 
2855=>X"0000010a0000010a0000010a0000010a", 2856=>X"0000010a0000010a0000010a0000010a", 2857=>X"0000010900000109000001090000010a", 2858=>X"00000109000001090000010900000109", 2859=>X"00000109000001090000010900000109", 
2860=>X"00000109000001090000010900000109", 2861=>X"00000108000001080000010800000108", 2862=>X"00000108000001080000010800000108", 2863=>X"00000108000001080000010800000108", 2864=>X"00000107000001080000010800000108", 
2865=>X"00000107000001070000010700000107", 2866=>X"00000107000001070000010700000107", 2867=>X"00000107000001070000010700000107", 2868=>X"00000106000001060000010700000107", 2869=>X"00000106000001060000010600000106", 
2870=>X"00000106000001060000010600000106", 2871=>X"00000106000001060000010600000106", 2872=>X"00000105000001050000010500000106", 2873=>X"00000105000001050000010500000105", 2874=>X"00000105000001050000010500000105", 
2875=>X"00000105000001050000010500000105", 2876=>X"00000104000001040000010400000105", 2877=>X"00000104000001040000010400000104", 2878=>X"00000104000001040000010400000104", 2879=>X"00000104000001040000010400000104", 
2880=>X"00000103000001030000010300000103", 2881=>X"00000103000001030000010300000103", 2882=>X"00000103000001030000010300000103", 2883=>X"00000103000001030000010300000103", 2884=>X"00000102000001020000010200000102", 
2885=>X"00000102000001020000010200000102", 2886=>X"00000102000001020000010200000102", 2887=>X"00000102000001020000010200000102", 2888=>X"00000101000001010000010100000101", 2889=>X"00000101000001010000010100000101", 
2890=>X"00000101000001010000010100000101", 2891=>X"00000101000001010000010100000101", 2892=>X"00000100000001000000010000000100", 2893=>X"00000100000001000000010000000100", 2894=>X"00000100000001000000010000000100", 
2895=>X"00000100000001000000010000000100", 2896=>X"000000ff000000ff000000ff000000ff", 2897=>X"000000ff000000ff000000ff000000ff", 2898=>X"000000ff000000ff000000ff000000ff", 2899=>X"000000ff000000ff000000ff000000ff", 
2900=>X"000000fe000000fe000000fe000000fe", 2901=>X"000000fe000000fe000000fe000000fe", 2902=>X"000000fe000000fe000000fe000000fe", 2903=>X"000000fe000000fe000000fe000000fe", 2904=>X"000000fd000000fd000000fd000000fd", 
2905=>X"000000fd000000fd000000fd000000fd", 2906=>X"000000fd000000fd000000fd000000fd", 2907=>X"000000fd000000fd000000fd000000fd", 2908=>X"000000fc000000fc000000fc000000fc", 2909=>X"000000fc000000fc000000fc000000fc", 
2910=>X"000000fc000000fc000000fc000000fc", 2911=>X"000000fc000000fc000000fc000000fc", 2912=>X"000000fb000000fb000000fb000000fc", 2913=>X"000000fb000000fb000000fb000000fb", 2914=>X"000000fb000000fb000000fb000000fb", 
2915=>X"000000fb000000fb000000fb000000fb", 2916=>X"000000fa000000fa000000fa000000fb", 2917=>X"000000fa000000fa000000fa000000fa", 2918=>X"000000fa000000fa000000fa000000fa", 2919=>X"000000fa000000fa000000fa000000fa", 
2920=>X"000000f9000000f9000000fa000000fa", 2921=>X"000000f9000000f9000000f9000000f9", 2922=>X"000000f9000000f9000000f9000000f9", 2923=>X"000000f9000000f9000000f9000000f9", 2924=>X"000000f8000000f9000000f9000000f9", 
2925=>X"000000f8000000f8000000f8000000f8", 2926=>X"000000f8000000f8000000f8000000f8", 2927=>X"000000f8000000f8000000f8000000f8", 2928=>X"000000f8000000f8000000f8000000f8", 2929=>X"000000f7000000f7000000f7000000f7", 
2930=>X"000000f7000000f7000000f7000000f7", 2931=>X"000000f7000000f7000000f7000000f7", 2932=>X"000000f7000000f7000000f7000000f7", 2933=>X"000000f6000000f6000000f6000000f7", 2934=>X"000000f6000000f6000000f6000000f6", 
2935=>X"000000f6000000f6000000f6000000f6", 2936=>X"000000f6000000f6000000f6000000f6", 2937=>X"000000f5000000f6000000f6000000f6", 2938=>X"000000f5000000f5000000f5000000f5", 2939=>X"000000f5000000f5000000f5000000f5", 
2940=>X"000000f5000000f5000000f5000000f5", 2941=>X"000000f5000000f5000000f5000000f5", 2942=>X"000000f4000000f4000000f4000000f4", 2943=>X"000000f4000000f4000000f4000000f4", 2944=>X"000000f4000000f4000000f4000000f4", 
2945=>X"000000f4000000f4000000f4000000f4", 2946=>X"000000f3000000f3000000f4000000f4", 2947=>X"000000f3000000f3000000f3000000f3", 2948=>X"000000f3000000f3000000f3000000f3", 2949=>X"000000f3000000f3000000f3000000f3", 
2950=>X"000000f3000000f3000000f3000000f3", 2951=>X"000000f2000000f2000000f2000000f2", 2952=>X"000000f2000000f2000000f2000000f2", 2953=>X"000000f2000000f2000000f2000000f2", 2954=>X"000000f2000000f2000000f2000000f2", 
2955=>X"000000f1000000f1000000f1000000f2", 2956=>X"000000f1000000f1000000f1000000f1", 2957=>X"000000f1000000f1000000f1000000f1", 2958=>X"000000f1000000f1000000f1000000f1", 2959=>X"000000f0000000f1000000f1000000f1", 
2960=>X"000000f0000000f0000000f0000000f0", 2961=>X"000000f0000000f0000000f0000000f0", 2962=>X"000000f0000000f0000000f0000000f0", 2963=>X"000000f0000000f0000000f0000000f0", 2964=>X"000000ef000000ef000000f0000000f0", 
2965=>X"000000ef000000ef000000ef000000ef", 2966=>X"000000ef000000ef000000ef000000ef", 2967=>X"000000ef000000ef000000ef000000ef", 2968=>X"000000ef000000ef000000ef000000ef", 2969=>X"000000ee000000ee000000ee000000ee", 
2970=>X"000000ee000000ee000000ee000000ee", 2971=>X"000000ee000000ee000000ee000000ee", 2972=>X"000000ee000000ee000000ee000000ee", 2973=>X"000000ed000000ee000000ee000000ee", 2974=>X"000000ed000000ed000000ed000000ed", 
2975=>X"000000ed000000ed000000ed000000ed", 2976=>X"000000ed000000ed000000ed000000ed", 2977=>X"000000ed000000ed000000ed000000ed", 2978=>X"000000ec000000ec000000ec000000ed", 2979=>X"000000ec000000ec000000ec000000ec", 
2980=>X"000000ec000000ec000000ec000000ec", 2981=>X"000000ec000000ec000000ec000000ec", 2982=>X"000000ec000000ec000000ec000000ec", 2983=>X"000000eb000000eb000000eb000000eb", 2984=>X"000000eb000000eb000000eb000000eb", 
2985=>X"000000eb000000eb000000eb000000eb", 2986=>X"000000eb000000eb000000eb000000eb", 2987=>X"000000ea000000eb000000eb000000eb", 2988=>X"000000ea000000ea000000ea000000ea", 2989=>X"000000ea000000ea000000ea000000ea", 
2990=>X"000000ea000000ea000000ea000000ea", 2991=>X"000000ea000000ea000000ea000000ea", 2992=>X"000000e9000000e9000000ea000000ea", 2993=>X"000000e9000000e9000000e9000000e9", 2994=>X"000000e9000000e9000000e9000000e9", 
2995=>X"000000e9000000e9000000e9000000e9", 2996=>X"000000e9000000e9000000e9000000e9", 2997=>X"000000e8000000e8000000e9000000e9", 2998=>X"000000e8000000e8000000e8000000e8", 2999=>X"000000e8000000e8000000e8000000e8", 
3000=>X"000000e8000000e8000000e8000000e8", 3001=>X"000000e8000000e8000000e8000000e8", 3002=>X"000000e7000000e7000000e7000000e8", 3003=>X"000000e7000000e7000000e7000000e7", 3004=>X"000000e7000000e7000000e7000000e7", 
3005=>X"000000e7000000e7000000e7000000e7", 3006=>X"000000e7000000e7000000e7000000e7", 3007=>X"000000e6000000e6000000e6000000e7", 3008=>X"000000e6000000e6000000e6000000e6", 3009=>X"000000e6000000e6000000e6000000e6", 
3010=>X"000000e6000000e6000000e6000000e6", 3011=>X"000000e6000000e6000000e6000000e6", 3012=>X"000000e5000000e5000000e5000000e5", 3013=>X"000000e5000000e5000000e5000000e5", 3014=>X"000000e5000000e5000000e5000000e5", 
3015=>X"000000e5000000e5000000e5000000e5", 3016=>X"000000e5000000e5000000e5000000e5", 3017=>X"000000e4000000e4000000e4000000e4", 3018=>X"000000e4000000e4000000e4000000e4", 3019=>X"000000e4000000e4000000e4000000e4", 
3020=>X"000000e4000000e4000000e4000000e4", 3021=>X"000000e4000000e4000000e4000000e4", 3022=>X"000000e3000000e3000000e3000000e4", 3023=>X"000000e3000000e3000000e3000000e3", 3024=>X"000000e3000000e3000000e3000000e3", 
3025=>X"000000e3000000e3000000e3000000e3", 3026=>X"000000e3000000e3000000e3000000e3", 3027=>X"000000e2000000e2000000e2000000e3", 3028=>X"000000e2000000e2000000e2000000e2", 3029=>X"000000e2000000e2000000e2000000e2", 
3030=>X"000000e2000000e2000000e2000000e2", 3031=>X"000000e2000000e2000000e2000000e2", 3032=>X"000000e1000000e1000000e2000000e2", 3033=>X"000000e1000000e1000000e1000000e1", 3034=>X"000000e1000000e1000000e1000000e1", 
3035=>X"000000e1000000e1000000e1000000e1", 3036=>X"000000e1000000e1000000e1000000e1", 3037=>X"000000e0000000e0000000e1000000e1", 3038=>X"000000e0000000e0000000e0000000e0", 3039=>X"000000e0000000e0000000e0000000e0", 
3040=>X"000000e0000000e0000000e0000000e0", 3041=>X"000000e0000000e0000000e0000000e0", 3042=>X"000000df000000e0000000e0000000e0", 3043=>X"000000df000000df000000df000000df", 3044=>X"000000df000000df000000df000000df", 
3045=>X"000000df000000df000000df000000df", 3046=>X"000000df000000df000000df000000df", 3047=>X"000000df000000df000000df000000df", 3048=>X"000000de000000de000000de000000de", 3049=>X"000000de000000de000000de000000de", 
3050=>X"000000de000000de000000de000000de", 3051=>X"000000de000000de000000de000000de", 3052=>X"000000de000000de000000de000000de", 3053=>X"000000dd000000dd000000dd000000de", 3054=>X"000000dd000000dd000000dd000000dd", 
3055=>X"000000dd000000dd000000dd000000dd", 3056=>X"000000dd000000dd000000dd000000dd", 3057=>X"000000dd000000dd000000dd000000dd", 3058=>X"000000dc000000dd000000dd000000dd", 3059=>X"000000dc000000dc000000dc000000dc", 
3060=>X"000000dc000000dc000000dc000000dc", 3061=>X"000000dc000000dc000000dc000000dc", 3062=>X"000000dc000000dc000000dc000000dc", 3063=>X"000000dc000000dc000000dc000000dc", 3064=>X"000000db000000db000000db000000dc", 
3065=>X"000000db000000db000000db000000db", 3066=>X"000000db000000db000000db000000db", 3067=>X"000000db000000db000000db000000db", 3068=>X"000000db000000db000000db000000db", 3069=>X"000000da000000da000000db000000db", 
3070=>X"000000da000000da000000da000000da", 3071=>X"000000da000000da000000da000000da", 3072=>X"000000da000000da000000da000000da", 3073=>X"000000da000000da000000da000000da", 3074=>X"000000da000000da000000da000000da", 
3075=>X"000000d9000000d9000000d9000000da", 3076=>X"000000d9000000d9000000d9000000d9", 3077=>X"000000d9000000d9000000d9000000d9", 3078=>X"000000d9000000d9000000d9000000d9", 3079=>X"000000d9000000d9000000d9000000d9", 
3080=>X"000000d8000000d9000000d9000000d9", 3081=>X"000000d8000000d8000000d8000000d8", 3082=>X"000000d8000000d8000000d8000000d8", 3083=>X"000000d8000000d8000000d8000000d8", 3084=>X"000000d8000000d8000000d8000000d8", 
3085=>X"000000d8000000d8000000d8000000d8", 3086=>X"000000d7000000d7000000d7000000d8", 3087=>X"000000d7000000d7000000d7000000d7", 3088=>X"000000d7000000d7000000d7000000d7", 3089=>X"000000d7000000d7000000d7000000d7", 
3090=>X"000000d7000000d7000000d7000000d7", 3091=>X"000000d7000000d7000000d7000000d7", 3092=>X"000000d6000000d6000000d6000000d6", 3093=>X"000000d6000000d6000000d6000000d6", 3094=>X"000000d6000000d6000000d6000000d6", 
3095=>X"000000d6000000d6000000d6000000d6", 3096=>X"000000d6000000d6000000d6000000d6", 3097=>X"000000d5000000d6000000d6000000d6", 3098=>X"000000d5000000d5000000d5000000d5", 3099=>X"000000d5000000d5000000d5000000d5", 
3100=>X"000000d5000000d5000000d5000000d5", 3101=>X"000000d5000000d5000000d5000000d5", 3102=>X"000000d5000000d5000000d5000000d5", 3103=>X"000000d4000000d4000000d5000000d5", 3104=>X"000000d4000000d4000000d4000000d4", 
3105=>X"000000d4000000d4000000d4000000d4", 3106=>X"000000d4000000d4000000d4000000d4", 3107=>X"000000d4000000d4000000d4000000d4", 3108=>X"000000d4000000d4000000d4000000d4", 3109=>X"000000d3000000d3000000d3000000d4", 
3110=>X"000000d3000000d3000000d3000000d3", 3111=>X"000000d3000000d3000000d3000000d3", 3112=>X"000000d3000000d3000000d3000000d3", 3113=>X"000000d3000000d3000000d3000000d3", 3114=>X"000000d3000000d3000000d3000000d3", 
3115=>X"000000d2000000d2000000d2000000d3", 3116=>X"000000d2000000d2000000d2000000d2", 3117=>X"000000d2000000d2000000d2000000d2", 3118=>X"000000d2000000d2000000d2000000d2", 3119=>X"000000d2000000d2000000d2000000d2", 
3120=>X"000000d2000000d2000000d2000000d2", 3121=>X"000000d1000000d1000000d1000000d2", 3122=>X"000000d1000000d1000000d1000000d1", 3123=>X"000000d1000000d1000000d1000000d1", 3124=>X"000000d1000000d1000000d1000000d1", 
3125=>X"000000d1000000d1000000d1000000d1", 3126=>X"000000d1000000d1000000d1000000d1", 3127=>X"000000d0000000d0000000d0000000d1", 3128=>X"000000d0000000d0000000d0000000d0", 3129=>X"000000d0000000d0000000d0000000d0", 
3130=>X"000000d0000000d0000000d0000000d0", 3131=>X"000000d0000000d0000000d0000000d0", 3132=>X"000000d0000000d0000000d0000000d0", 3133=>X"000000cf000000cf000000cf000000d0", 3134=>X"000000cf000000cf000000cf000000cf", 
3135=>X"000000cf000000cf000000cf000000cf", 3136=>X"000000cf000000cf000000cf000000cf", 3137=>X"000000cf000000cf000000cf000000cf", 3138=>X"000000cf000000cf000000cf000000cf", 3139=>X"000000ce000000ce000000ce000000cf", 
3140=>X"000000ce000000ce000000ce000000ce", 3141=>X"000000ce000000ce000000ce000000ce", 3142=>X"000000ce000000ce000000ce000000ce", 3143=>X"000000ce000000ce000000ce000000ce", 3144=>X"000000ce000000ce000000ce000000ce", 
3145=>X"000000cd000000cd000000ce000000ce", 3146=>X"000000cd000000cd000000cd000000cd", 3147=>X"000000cd000000cd000000cd000000cd", 3148=>X"000000cd000000cd000000cd000000cd", 3149=>X"000000cd000000cd000000cd000000cd", 
3150=>X"000000cd000000cd000000cd000000cd", 3151=>X"000000cc000000cd000000cd000000cd", 3152=>X"000000cc000000cc000000cc000000cc", 3153=>X"000000cc000000cc000000cc000000cc", 3154=>X"000000cc000000cc000000cc000000cc", 
3155=>X"000000cc000000cc000000cc000000cc", 3156=>X"000000cc000000cc000000cc000000cc", 3157=>X"000000cc000000cc000000cc000000cc", 3158=>X"000000cb000000cb000000cb000000cb", 3159=>X"000000cb000000cb000000cb000000cb", 
3160=>X"000000cb000000cb000000cb000000cb", 3161=>X"000000cb000000cb000000cb000000cb", 3162=>X"000000cb000000cb000000cb000000cb", 3163=>X"000000cb000000cb000000cb000000cb", 3164=>X"000000ca000000ca000000cb000000cb", 
3165=>X"000000ca000000ca000000ca000000ca", 3166=>X"000000ca000000ca000000ca000000ca", 3167=>X"000000ca000000ca000000ca000000ca", 3168=>X"000000ca000000ca000000ca000000ca", 3169=>X"000000ca000000ca000000ca000000ca", 
3170=>X"000000c9000000ca000000ca000000ca", 3171=>X"000000c9000000c9000000c9000000c9", 3172=>X"000000c9000000c9000000c9000000c9", 3173=>X"000000c9000000c9000000c9000000c9", 3174=>X"000000c9000000c9000000c9000000c9", 
3175=>X"000000c9000000c9000000c9000000c9", 3176=>X"000000c9000000c9000000c9000000c9", 3177=>X"000000c8000000c8000000c8000000c9", 3178=>X"000000c8000000c8000000c8000000c8", 3179=>X"000000c8000000c8000000c8000000c8", 
3180=>X"000000c8000000c8000000c8000000c8", 3181=>X"000000c8000000c8000000c8000000c8", 3182=>X"000000c8000000c8000000c8000000c8", 3183=>X"000000c8000000c8000000c8000000c8", 3184=>X"000000c7000000c7000000c7000000c7", 
3185=>X"000000c7000000c7000000c7000000c7", 3186=>X"000000c7000000c7000000c7000000c7", 3187=>X"000000c7000000c7000000c7000000c7", 3188=>X"000000c7000000c7000000c7000000c7", 3189=>X"000000c7000000c7000000c7000000c7", 
3190=>X"000000c6000000c6000000c7000000c7", 3191=>X"000000c6000000c6000000c6000000c6", 3192=>X"000000c6000000c6000000c6000000c6", 3193=>X"000000c6000000c6000000c6000000c6", 3194=>X"000000c6000000c6000000c6000000c6", 
3195=>X"000000c6000000c6000000c6000000c6", 3196=>X"000000c6000000c6000000c6000000c6", 3197=>X"000000c5000000c5000000c5000000c6", 3198=>X"000000c5000000c5000000c5000000c5", 3199=>X"000000c5000000c5000000c5000000c5", 
3200=>X"000000c5000000c5000000c5000000c5", 3201=>X"000000c5000000c5000000c5000000c5", 3202=>X"000000c5000000c5000000c5000000c5", 3203=>X"000000c5000000c5000000c5000000c5", 3204=>X"000000c4000000c4000000c4000000c4", 
3205=>X"000000c4000000c4000000c4000000c4", 3206=>X"000000c4000000c4000000c4000000c4", 3207=>X"000000c4000000c4000000c4000000c4", 3208=>X"000000c4000000c4000000c4000000c4", 3209=>X"000000c4000000c4000000c4000000c4", 
3210=>X"000000c3000000c4000000c4000000c4", 3211=>X"000000c3000000c3000000c3000000c3", 3212=>X"000000c3000000c3000000c3000000c3", 3213=>X"000000c3000000c3000000c3000000c3", 3214=>X"000000c3000000c3000000c3000000c3", 
3215=>X"000000c3000000c3000000c3000000c3", 3216=>X"000000c3000000c3000000c3000000c3", 3217=>X"000000c2000000c3000000c3000000c3", 3218=>X"000000c2000000c2000000c2000000c2", 3219=>X"000000c2000000c2000000c2000000c2", 
3220=>X"000000c2000000c2000000c2000000c2", 3221=>X"000000c2000000c2000000c2000000c2", 3222=>X"000000c2000000c2000000c2000000c2", 3223=>X"000000c2000000c2000000c2000000c2", 3224=>X"000000c1000000c1000000c2000000c2", 
3225=>X"000000c1000000c1000000c1000000c1", 3226=>X"000000c1000000c1000000c1000000c1", 3227=>X"000000c1000000c1000000c1000000c1", 3228=>X"000000c1000000c1000000c1000000c1", 3229=>X"000000c1000000c1000000c1000000c1", 
3230=>X"000000c1000000c1000000c1000000c1", 3231=>X"000000c0000000c1000000c1000000c1", 3232=>X"000000c0000000c0000000c0000000c0", 3233=>X"000000c0000000c0000000c0000000c0", 3234=>X"000000c0000000c0000000c0000000c0", 
3235=>X"000000c0000000c0000000c0000000c0", 3236=>X"000000c0000000c0000000c0000000c0", 3237=>X"000000c0000000c0000000c0000000c0", 3238=>X"000000bf000000c0000000c0000000c0", 3239=>X"000000bf000000bf000000bf000000bf", 
3240=>X"000000bf000000bf000000bf000000bf", 3241=>X"000000bf000000bf000000bf000000bf", 3242=>X"000000bf000000bf000000bf000000bf", 3243=>X"000000bf000000bf000000bf000000bf", 3244=>X"000000bf000000bf000000bf000000bf", 
3245=>X"000000bf000000bf000000bf000000bf", 3246=>X"000000be000000be000000be000000be", 3247=>X"000000be000000be000000be000000be", 3248=>X"000000be000000be000000be000000be", 3249=>X"000000be000000be000000be000000be", 
3250=>X"000000be000000be000000be000000be", 3251=>X"000000be000000be000000be000000be", 3252=>X"000000be000000be000000be000000be", 3253=>X"000000bd000000bd000000bd000000be", 3254=>X"000000bd000000bd000000bd000000bd", 
3255=>X"000000bd000000bd000000bd000000bd", 3256=>X"000000bd000000bd000000bd000000bd", 3257=>X"000000bd000000bd000000bd000000bd", 3258=>X"000000bd000000bd000000bd000000bd", 3259=>X"000000bd000000bd000000bd000000bd", 
3260=>X"000000bc000000bc000000bd000000bd", 3261=>X"000000bc000000bc000000bc000000bc", 3262=>X"000000bc000000bc000000bc000000bc", 3263=>X"000000bc000000bc000000bc000000bc", 3264=>X"000000bc000000bc000000bc000000bc", 
3265=>X"000000bc000000bc000000bc000000bc", 3266=>X"000000bc000000bc000000bc000000bc", 3267=>X"000000bc000000bc000000bc000000bc", 3268=>X"000000bb000000bb000000bb000000bb", 3269=>X"000000bb000000bb000000bb000000bb", 
3270=>X"000000bb000000bb000000bb000000bb", 3271=>X"000000bb000000bb000000bb000000bb", 3272=>X"000000bb000000bb000000bb000000bb", 3273=>X"000000bb000000bb000000bb000000bb", 3274=>X"000000bb000000bb000000bb000000bb", 
3275=>X"000000ba000000ba000000bb000000bb", 3276=>X"000000ba000000ba000000ba000000ba", 3277=>X"000000ba000000ba000000ba000000ba", 3278=>X"000000ba000000ba000000ba000000ba", 3279=>X"000000ba000000ba000000ba000000ba", 
3280=>X"000000ba000000ba000000ba000000ba", 3281=>X"000000ba000000ba000000ba000000ba", 3282=>X"000000ba000000ba000000ba000000ba", 3283=>X"000000b9000000b9000000b9000000b9", 3284=>X"000000b9000000b9000000b9000000b9", 
3285=>X"000000b9000000b9000000b9000000b9", 3286=>X"000000b9000000b9000000b9000000b9", 3287=>X"000000b9000000b9000000b9000000b9", 3288=>X"000000b9000000b9000000b9000000b9", 3289=>X"000000b9000000b9000000b9000000b9", 
3290=>X"000000b8000000b9000000b9000000b9", 3291=>X"000000b8000000b8000000b8000000b8", 3292=>X"000000b8000000b8000000b8000000b8", 3293=>X"000000b8000000b8000000b8000000b8", 3294=>X"000000b8000000b8000000b8000000b8", 
3295=>X"000000b8000000b8000000b8000000b8", 3296=>X"000000b8000000b8000000b8000000b8", 3297=>X"000000b8000000b8000000b8000000b8", 3298=>X"000000b7000000b7000000b8000000b8", 3299=>X"000000b7000000b7000000b7000000b7", 
3300=>X"000000b7000000b7000000b7000000b7", 3301=>X"000000b7000000b7000000b7000000b7", 3302=>X"000000b7000000b7000000b7000000b7", 3303=>X"000000b7000000b7000000b7000000b7", 3304=>X"000000b7000000b7000000b7000000b7", 
3305=>X"000000b7000000b7000000b7000000b7", 3306=>X"000000b6000000b6000000b6000000b7", 3307=>X"000000b6000000b6000000b6000000b6", 3308=>X"000000b6000000b6000000b6000000b6", 3309=>X"000000b6000000b6000000b6000000b6", 
3310=>X"000000b6000000b6000000b6000000b6", 3311=>X"000000b6000000b6000000b6000000b6", 3312=>X"000000b6000000b6000000b6000000b6", 3313=>X"000000b6000000b6000000b6000000b6", 3314=>X"000000b5000000b5000000b5000000b6", 
3315=>X"000000b5000000b5000000b5000000b5", 3316=>X"000000b5000000b5000000b5000000b5", 3317=>X"000000b5000000b5000000b5000000b5", 3318=>X"000000b5000000b5000000b5000000b5", 3319=>X"000000b5000000b5000000b5000000b5", 
3320=>X"000000b5000000b5000000b5000000b5", 3321=>X"000000b5000000b5000000b5000000b5", 3322=>X"000000b4000000b4000000b4000000b5", 3323=>X"000000b4000000b4000000b4000000b4", 3324=>X"000000b4000000b4000000b4000000b4", 
3325=>X"000000b4000000b4000000b4000000b4", 3326=>X"000000b4000000b4000000b4000000b4", 3327=>X"000000b4000000b4000000b4000000b4", 3328=>X"000000b4000000b4000000b4000000b4", 3329=>X"000000b4000000b4000000b4000000b4", 
3330=>X"000000b3000000b3000000b3000000b4", 3331=>X"000000b3000000b3000000b3000000b3", 3332=>X"000000b3000000b3000000b3000000b3", 3333=>X"000000b3000000b3000000b3000000b3", 3334=>X"000000b3000000b3000000b3000000b3", 
3335=>X"000000b3000000b3000000b3000000b3", 3336=>X"000000b3000000b3000000b3000000b3", 3337=>X"000000b3000000b3000000b3000000b3", 3338=>X"000000b2000000b2000000b3000000b3", 3339=>X"000000b2000000b2000000b2000000b2", 
3340=>X"000000b2000000b2000000b2000000b2", 3341=>X"000000b2000000b2000000b2000000b2", 3342=>X"000000b2000000b2000000b2000000b2", 3343=>X"000000b2000000b2000000b2000000b2", 3344=>X"000000b2000000b2000000b2000000b2", 
3345=>X"000000b2000000b2000000b2000000b2", 3346=>X"000000b1000000b2000000b2000000b2", 3347=>X"000000b1000000b1000000b1000000b1", 3348=>X"000000b1000000b1000000b1000000b1", 3349=>X"000000b1000000b1000000b1000000b1", 
3350=>X"000000b1000000b1000000b1000000b1", 3351=>X"000000b1000000b1000000b1000000b1", 3352=>X"000000b1000000b1000000b1000000b1", 3353=>X"000000b1000000b1000000b1000000b1", 3354=>X"000000b1000000b1000000b1000000b1", 
3355=>X"000000b0000000b0000000b0000000b0", 3356=>X"000000b0000000b0000000b0000000b0", 3357=>X"000000b0000000b0000000b0000000b0", 3358=>X"000000b0000000b0000000b0000000b0", 3359=>X"000000b0000000b0000000b0000000b0", 
3360=>X"000000b0000000b0000000b0000000b0", 3361=>X"000000b0000000b0000000b0000000b0", 3362=>X"000000b0000000b0000000b0000000b0", 3363=>X"000000af000000af000000b0000000b0", 3364=>X"000000af000000af000000af000000af", 
3365=>X"000000af000000af000000af000000af", 3366=>X"000000af000000af000000af000000af", 3367=>X"000000af000000af000000af000000af", 3368=>X"000000af000000af000000af000000af", 3369=>X"000000af000000af000000af000000af", 
3370=>X"000000af000000af000000af000000af", 3371=>X"000000af000000af000000af000000af", 3372=>X"000000ae000000ae000000ae000000af", 3373=>X"000000ae000000ae000000ae000000ae", 3374=>X"000000ae000000ae000000ae000000ae", 
3375=>X"000000ae000000ae000000ae000000ae", 3376=>X"000000ae000000ae000000ae000000ae", 3377=>X"000000ae000000ae000000ae000000ae", 3378=>X"000000ae000000ae000000ae000000ae", 3379=>X"000000ae000000ae000000ae000000ae", 
3380=>X"000000ad000000ae000000ae000000ae", 3381=>X"000000ad000000ad000000ad000000ad", 3382=>X"000000ad000000ad000000ad000000ad", 3383=>X"000000ad000000ad000000ad000000ad", 3384=>X"000000ad000000ad000000ad000000ad", 
3385=>X"000000ad000000ad000000ad000000ad", 3386=>X"000000ad000000ad000000ad000000ad", 3387=>X"000000ad000000ad000000ad000000ad", 3388=>X"000000ad000000ad000000ad000000ad", 3389=>X"000000ac000000ac000000ad000000ad", 
3390=>X"000000ac000000ac000000ac000000ac", 3391=>X"000000ac000000ac000000ac000000ac", 3392=>X"000000ac000000ac000000ac000000ac", 3393=>X"000000ac000000ac000000ac000000ac", 3394=>X"000000ac000000ac000000ac000000ac", 
3395=>X"000000ac000000ac000000ac000000ac", 3396=>X"000000ac000000ac000000ac000000ac", 3397=>X"000000ac000000ac000000ac000000ac", 3398=>X"000000ab000000ab000000ac000000ac", 3399=>X"000000ab000000ab000000ab000000ab", 
3400=>X"000000ab000000ab000000ab000000ab", 3401=>X"000000ab000000ab000000ab000000ab", 3402=>X"000000ab000000ab000000ab000000ab", 3403=>X"000000ab000000ab000000ab000000ab", 3404=>X"000000ab000000ab000000ab000000ab", 
3405=>X"000000ab000000ab000000ab000000ab", 3406=>X"000000ab000000ab000000ab000000ab", 3407=>X"000000aa000000aa000000ab000000ab", 3408=>X"000000aa000000aa000000aa000000aa", 3409=>X"000000aa000000aa000000aa000000aa", 
3410=>X"000000aa000000aa000000aa000000aa", 3411=>X"000000aa000000aa000000aa000000aa", 3412=>X"000000aa000000aa000000aa000000aa", 3413=>X"000000aa000000aa000000aa000000aa", 3414=>X"000000aa000000aa000000aa000000aa", 
3415=>X"000000aa000000aa000000aa000000aa", 3416=>X"000000a9000000a9000000aa000000aa", 3417=>X"000000a9000000a9000000a9000000a9", 3418=>X"000000a9000000a9000000a9000000a9", 3419=>X"000000a9000000a9000000a9000000a9", 
3420=>X"000000a9000000a9000000a9000000a9", 3421=>X"000000a9000000a9000000a9000000a9", 3422=>X"000000a9000000a9000000a9000000a9", 3423=>X"000000a9000000a9000000a9000000a9", 3424=>X"000000a9000000a9000000a9000000a9", 
3425=>X"000000a8000000a9000000a9000000a9", 3426=>X"000000a8000000a8000000a8000000a8", 3427=>X"000000a8000000a8000000a8000000a8", 3428=>X"000000a8000000a8000000a8000000a8", 3429=>X"000000a8000000a8000000a8000000a8", 
3430=>X"000000a8000000a8000000a8000000a8", 3431=>X"000000a8000000a8000000a8000000a8", 3432=>X"000000a8000000a8000000a8000000a8", 3433=>X"000000a8000000a8000000a8000000a8", 3434=>X"000000a8000000a8000000a8000000a8", 
3435=>X"000000a7000000a7000000a7000000a7", 3436=>X"000000a7000000a7000000a7000000a7", 3437=>X"000000a7000000a7000000a7000000a7", 3438=>X"000000a7000000a7000000a7000000a7", 3439=>X"000000a7000000a7000000a7000000a7", 
3440=>X"000000a7000000a7000000a7000000a7", 3441=>X"000000a7000000a7000000a7000000a7", 3442=>X"000000a7000000a7000000a7000000a7", 3443=>X"000000a7000000a7000000a7000000a7", 3444=>X"000000a6000000a6000000a6000000a7", 
3445=>X"000000a6000000a6000000a6000000a6", 3446=>X"000000a6000000a6000000a6000000a6", 3447=>X"000000a6000000a6000000a6000000a6", 3448=>X"000000a6000000a6000000a6000000a6", 3449=>X"000000a6000000a6000000a6000000a6", 
3450=>X"000000a6000000a6000000a6000000a6", 3451=>X"000000a6000000a6000000a6000000a6", 3452=>X"000000a6000000a6000000a6000000a6", 3453=>X"000000a5000000a6000000a6000000a6", 3454=>X"000000a5000000a5000000a5000000a5", 
3455=>X"000000a5000000a5000000a5000000a5", 3456=>X"000000a5000000a5000000a5000000a5", 3457=>X"000000a5000000a5000000a5000000a5", 3458=>X"000000a5000000a5000000a5000000a5", 3459=>X"000000a5000000a5000000a5000000a5", 
3460=>X"000000a5000000a5000000a5000000a5", 3461=>X"000000a5000000a5000000a5000000a5", 3462=>X"000000a5000000a5000000a5000000a5", 3463=>X"000000a4000000a4000000a5000000a5", 3464=>X"000000a4000000a4000000a4000000a4", 
3465=>X"000000a4000000a4000000a4000000a4", 3466=>X"000000a4000000a4000000a4000000a4", 3467=>X"000000a4000000a4000000a4000000a4", 3468=>X"000000a4000000a4000000a4000000a4", 3469=>X"000000a4000000a4000000a4000000a4", 
3470=>X"000000a4000000a4000000a4000000a4", 3471=>X"000000a4000000a4000000a4000000a4", 3472=>X"000000a4000000a4000000a4000000a4", 3473=>X"000000a3000000a3000000a3000000a4", 3474=>X"000000a3000000a3000000a3000000a3", 
3475=>X"000000a3000000a3000000a3000000a3", 3476=>X"000000a3000000a3000000a3000000a3", 3477=>X"000000a3000000a3000000a3000000a3", 3478=>X"000000a3000000a3000000a3000000a3", 3479=>X"000000a3000000a3000000a3000000a3", 
3480=>X"000000a3000000a3000000a3000000a3", 3481=>X"000000a3000000a3000000a3000000a3", 3482=>X"000000a3000000a3000000a3000000a3", 3483=>X"000000a2000000a2000000a2000000a2", 3484=>X"000000a2000000a2000000a2000000a2", 
3485=>X"000000a2000000a2000000a2000000a2", 3486=>X"000000a2000000a2000000a2000000a2", 3487=>X"000000a2000000a2000000a2000000a2", 3488=>X"000000a2000000a2000000a2000000a2", 3489=>X"000000a2000000a2000000a2000000a2", 
3490=>X"000000a2000000a2000000a2000000a2", 3491=>X"000000a2000000a2000000a2000000a2", 3492=>X"000000a2000000a2000000a2000000a2", 3493=>X"000000a1000000a1000000a1000000a1", 3494=>X"000000a1000000a1000000a1000000a1", 
3495=>X"000000a1000000a1000000a1000000a1", 3496=>X"000000a1000000a1000000a1000000a1", 3497=>X"000000a1000000a1000000a1000000a1", 3498=>X"000000a1000000a1000000a1000000a1", 3499=>X"000000a1000000a1000000a1000000a1", 
3500=>X"000000a1000000a1000000a1000000a1", 3501=>X"000000a1000000a1000000a1000000a1", 3502=>X"000000a1000000a1000000a1000000a1", 3503=>X"000000a0000000a0000000a0000000a1", 3504=>X"000000a0000000a0000000a0000000a0", 
3505=>X"000000a0000000a0000000a0000000a0", 3506=>X"000000a0000000a0000000a0000000a0", 3507=>X"000000a0000000a0000000a0000000a0", 3508=>X"000000a0000000a0000000a0000000a0", 3509=>X"000000a0000000a0000000a0000000a0", 
3510=>X"000000a0000000a0000000a0000000a0", 3511=>X"000000a0000000a0000000a0000000a0", 3512=>X"000000a0000000a0000000a0000000a0", 3513=>X"0000009f0000009f000000a0000000a0", 3514=>X"0000009f0000009f0000009f0000009f", 
3515=>X"0000009f0000009f0000009f0000009f", 3516=>X"0000009f0000009f0000009f0000009f", 3517=>X"0000009f0000009f0000009f0000009f", 3518=>X"0000009f0000009f0000009f0000009f", 3519=>X"0000009f0000009f0000009f0000009f", 
3520=>X"0000009f0000009f0000009f0000009f", 3521=>X"0000009f0000009f0000009f0000009f", 3522=>X"0000009f0000009f0000009f0000009f", 3523=>X"0000009e0000009f0000009f0000009f", 3524=>X"0000009e0000009e0000009e0000009e", 
3525=>X"0000009e0000009e0000009e0000009e", 3526=>X"0000009e0000009e0000009e0000009e", 3527=>X"0000009e0000009e0000009e0000009e", 3528=>X"0000009e0000009e0000009e0000009e", 3529=>X"0000009e0000009e0000009e0000009e", 
3530=>X"0000009e0000009e0000009e0000009e", 3531=>X"0000009e0000009e0000009e0000009e", 3532=>X"0000009e0000009e0000009e0000009e", 3533=>X"0000009e0000009e0000009e0000009e", 3534=>X"0000009d0000009d0000009d0000009e", 
3535=>X"0000009d0000009d0000009d0000009d", 3536=>X"0000009d0000009d0000009d0000009d", 3537=>X"0000009d0000009d0000009d0000009d", 3538=>X"0000009d0000009d0000009d0000009d", 3539=>X"0000009d0000009d0000009d0000009d", 
3540=>X"0000009d0000009d0000009d0000009d", 3541=>X"0000009d0000009d0000009d0000009d", 3542=>X"0000009d0000009d0000009d0000009d", 3543=>X"0000009d0000009d0000009d0000009d", 3544=>X"0000009d0000009d0000009d0000009d", 
3545=>X"0000009c0000009c0000009c0000009c", 3546=>X"0000009c0000009c0000009c0000009c", 3547=>X"0000009c0000009c0000009c0000009c", 3548=>X"0000009c0000009c0000009c0000009c", 3549=>X"0000009c0000009c0000009c0000009c", 
3550=>X"0000009c0000009c0000009c0000009c", 3551=>X"0000009c0000009c0000009c0000009c", 3552=>X"0000009c0000009c0000009c0000009c", 3553=>X"0000009c0000009c0000009c0000009c", 3554=>X"0000009c0000009c0000009c0000009c", 
3555=>X"0000009b0000009c0000009c0000009c", 3556=>X"0000009b0000009b0000009b0000009b", 3557=>X"0000009b0000009b0000009b0000009b", 3558=>X"0000009b0000009b0000009b0000009b", 3559=>X"0000009b0000009b0000009b0000009b", 
3560=>X"0000009b0000009b0000009b0000009b", 3561=>X"0000009b0000009b0000009b0000009b", 3562=>X"0000009b0000009b0000009b0000009b", 3563=>X"0000009b0000009b0000009b0000009b", 3564=>X"0000009b0000009b0000009b0000009b", 
3565=>X"0000009b0000009b0000009b0000009b", 3566=>X"0000009a0000009a0000009b0000009b", 3567=>X"0000009a0000009a0000009a0000009a", 3568=>X"0000009a0000009a0000009a0000009a", 3569=>X"0000009a0000009a0000009a0000009a", 
3570=>X"0000009a0000009a0000009a0000009a", 3571=>X"0000009a0000009a0000009a0000009a", 3572=>X"0000009a0000009a0000009a0000009a", 3573=>X"0000009a0000009a0000009a0000009a", 3574=>X"0000009a0000009a0000009a0000009a", 
3575=>X"0000009a0000009a0000009a0000009a", 3576=>X"0000009a0000009a0000009a0000009a", 3577=>X"000000990000009a0000009a0000009a", 3578=>X"00000099000000990000009900000099", 3579=>X"00000099000000990000009900000099", 
3580=>X"00000099000000990000009900000099", 3581=>X"00000099000000990000009900000099", 3582=>X"00000099000000990000009900000099", 3583=>X"00000099000000990000009900000099", 3584=>X"00000099000000990000009900000099", 
3585=>X"00000099000000990000009900000099", 3586=>X"00000099000000990000009900000099", 3587=>X"00000099000000990000009900000099", 3588=>X"00000098000000990000009900000099", 3589=>X"00000098000000980000009800000098", 
3590=>X"00000098000000980000009800000098", 3591=>X"00000098000000980000009800000098", 3592=>X"00000098000000980000009800000098", 3593=>X"00000098000000980000009800000098", 3594=>X"00000098000000980000009800000098", 
3595=>X"00000098000000980000009800000098", 3596=>X"00000098000000980000009800000098", 3597=>X"00000098000000980000009800000098", 3598=>X"00000098000000980000009800000098", 3599=>X"00000098000000980000009800000098", 
3600=>X"00000097000000970000009700000098", 3601=>X"00000097000000970000009700000097", 3602=>X"00000097000000970000009700000097", 3603=>X"00000097000000970000009700000097", 3604=>X"00000097000000970000009700000097", 
3605=>X"00000097000000970000009700000097", 3606=>X"00000097000000970000009700000097", 3607=>X"00000097000000970000009700000097", 3608=>X"00000097000000970000009700000097", 3609=>X"00000097000000970000009700000097", 
3610=>X"00000097000000970000009700000097", 3611=>X"00000096000000970000009700000097", 3612=>X"00000096000000960000009600000096", 3613=>X"00000096000000960000009600000096", 3614=>X"00000096000000960000009600000096", 
3615=>X"00000096000000960000009600000096", 3616=>X"00000096000000960000009600000096", 3617=>X"00000096000000960000009600000096", 3618=>X"00000096000000960000009600000096", 3619=>X"00000096000000960000009600000096", 
3620=>X"00000096000000960000009600000096", 3621=>X"00000096000000960000009600000096", 3622=>X"00000096000000960000009600000096", 3623=>X"00000095000000950000009500000096", 3624=>X"00000095000000950000009500000095", 
3625=>X"00000095000000950000009500000095", 3626=>X"00000095000000950000009500000095", 3627=>X"00000095000000950000009500000095", 3628=>X"00000095000000950000009500000095", 3629=>X"00000095000000950000009500000095", 
3630=>X"00000095000000950000009500000095", 3631=>X"00000095000000950000009500000095", 3632=>X"00000095000000950000009500000095", 3633=>X"00000095000000950000009500000095", 3634=>X"00000095000000950000009500000095", 
3635=>X"00000094000000940000009400000095", 3636=>X"00000094000000940000009400000094", 3637=>X"00000094000000940000009400000094", 3638=>X"00000094000000940000009400000094", 3639=>X"00000094000000940000009400000094", 
3640=>X"00000094000000940000009400000094", 3641=>X"00000094000000940000009400000094", 3642=>X"00000094000000940000009400000094", 3643=>X"00000094000000940000009400000094", 3644=>X"00000094000000940000009400000094", 
3645=>X"00000094000000940000009400000094", 3646=>X"00000094000000940000009400000094", 3647=>X"00000093000000930000009300000093", 3648=>X"00000093000000930000009300000093", 3649=>X"00000093000000930000009300000093", 
3650=>X"00000093000000930000009300000093", 3651=>X"00000093000000930000009300000093", 3652=>X"00000093000000930000009300000093", 3653=>X"00000093000000930000009300000093", 3654=>X"00000093000000930000009300000093", 
3655=>X"00000093000000930000009300000093", 3656=>X"00000093000000930000009300000093", 3657=>X"00000093000000930000009300000093", 3658=>X"00000093000000930000009300000093", 3659=>X"00000092000000920000009200000093", 
3660=>X"00000092000000920000009200000092", 3661=>X"00000092000000920000009200000092", 3662=>X"00000092000000920000009200000092", 3663=>X"00000092000000920000009200000092", 3664=>X"00000092000000920000009200000092", 
3665=>X"00000092000000920000009200000092", 3666=>X"00000092000000920000009200000092", 3667=>X"00000092000000920000009200000092", 3668=>X"00000092000000920000009200000092", 3669=>X"00000092000000920000009200000092", 
3670=>X"00000092000000920000009200000092", 3671=>X"00000091000000910000009200000092", 3672=>X"00000091000000910000009100000091", 3673=>X"00000091000000910000009100000091", 3674=>X"00000091000000910000009100000091", 
3675=>X"00000091000000910000009100000091", 3676=>X"00000091000000910000009100000091", 3677=>X"00000091000000910000009100000091", 3678=>X"00000091000000910000009100000091", 3679=>X"00000091000000910000009100000091", 
3680=>X"00000091000000910000009100000091", 3681=>X"00000091000000910000009100000091", 3682=>X"00000091000000910000009100000091", 3683=>X"00000091000000910000009100000091", 3684=>X"00000090000000900000009000000090", 
3685=>X"00000090000000900000009000000090", 3686=>X"00000090000000900000009000000090", 3687=>X"00000090000000900000009000000090", 3688=>X"00000090000000900000009000000090", 3689=>X"00000090000000900000009000000090", 
3690=>X"00000090000000900000009000000090", 3691=>X"00000090000000900000009000000090", 3692=>X"00000090000000900000009000000090", 3693=>X"00000090000000900000009000000090", 3694=>X"00000090000000900000009000000090", 
3695=>X"00000090000000900000009000000090", 3696=>X"0000008f000000900000009000000090", 3697=>X"0000008f0000008f0000008f0000008f", 3698=>X"0000008f0000008f0000008f0000008f", 3699=>X"0000008f0000008f0000008f0000008f", 
3700=>X"0000008f0000008f0000008f0000008f", 3701=>X"0000008f0000008f0000008f0000008f", 3702=>X"0000008f0000008f0000008f0000008f", 3703=>X"0000008f0000008f0000008f0000008f", 3704=>X"0000008f0000008f0000008f0000008f", 
3705=>X"0000008f0000008f0000008f0000008f", 3706=>X"0000008f0000008f0000008f0000008f", 3707=>X"0000008f0000008f0000008f0000008f", 3708=>X"0000008f0000008f0000008f0000008f", 3709=>X"0000008e0000008e0000008f0000008f", 
3710=>X"0000008e0000008e0000008e0000008e", 3711=>X"0000008e0000008e0000008e0000008e", 3712=>X"0000008e0000008e0000008e0000008e", 3713=>X"0000008e0000008e0000008e0000008e", 3714=>X"0000008e0000008e0000008e0000008e", 
3715=>X"0000008e0000008e0000008e0000008e", 3716=>X"0000008e0000008e0000008e0000008e", 3717=>X"0000008e0000008e0000008e0000008e", 3718=>X"0000008e0000008e0000008e0000008e", 3719=>X"0000008e0000008e0000008e0000008e", 
3720=>X"0000008e0000008e0000008e0000008e", 3721=>X"0000008e0000008e0000008e0000008e", 3722=>X"0000008d0000008d0000008e0000008e", 3723=>X"0000008d0000008d0000008d0000008d", 3724=>X"0000008d0000008d0000008d0000008d", 
3725=>X"0000008d0000008d0000008d0000008d", 3726=>X"0000008d0000008d0000008d0000008d", 3727=>X"0000008d0000008d0000008d0000008d", 3728=>X"0000008d0000008d0000008d0000008d", 3729=>X"0000008d0000008d0000008d0000008d", 
3730=>X"0000008d0000008d0000008d0000008d", 3731=>X"0000008d0000008d0000008d0000008d", 3732=>X"0000008d0000008d0000008d0000008d", 3733=>X"0000008d0000008d0000008d0000008d", 3734=>X"0000008d0000008d0000008d0000008d", 
3735=>X"0000008c0000008d0000008d0000008d", 3736=>X"0000008c0000008c0000008c0000008c", 3737=>X"0000008c0000008c0000008c0000008c", 3738=>X"0000008c0000008c0000008c0000008c", 3739=>X"0000008c0000008c0000008c0000008c", 
3740=>X"0000008c0000008c0000008c0000008c", 3741=>X"0000008c0000008c0000008c0000008c", 3742=>X"0000008c0000008c0000008c0000008c", 3743=>X"0000008c0000008c0000008c0000008c", 3744=>X"0000008c0000008c0000008c0000008c", 
3745=>X"0000008c0000008c0000008c0000008c", 3746=>X"0000008c0000008c0000008c0000008c", 3747=>X"0000008c0000008c0000008c0000008c", 3748=>X"0000008c0000008c0000008c0000008c", 3749=>X"0000008b0000008b0000008b0000008b", 
3750=>X"0000008b0000008b0000008b0000008b", 3751=>X"0000008b0000008b0000008b0000008b", 3752=>X"0000008b0000008b0000008b0000008b", 3753=>X"0000008b0000008b0000008b0000008b", 3754=>X"0000008b0000008b0000008b0000008b", 
3755=>X"0000008b0000008b0000008b0000008b", 3756=>X"0000008b0000008b0000008b0000008b", 3757=>X"0000008b0000008b0000008b0000008b", 3758=>X"0000008b0000008b0000008b0000008b", 3759=>X"0000008b0000008b0000008b0000008b", 
3760=>X"0000008b0000008b0000008b0000008b", 3761=>X"0000008b0000008b0000008b0000008b", 3762=>X"0000008a0000008a0000008b0000008b", 3763=>X"0000008a0000008a0000008a0000008a", 3764=>X"0000008a0000008a0000008a0000008a", 
3765=>X"0000008a0000008a0000008a0000008a", 3766=>X"0000008a0000008a0000008a0000008a", 3767=>X"0000008a0000008a0000008a0000008a", 3768=>X"0000008a0000008a0000008a0000008a", 3769=>X"0000008a0000008a0000008a0000008a", 
3770=>X"0000008a0000008a0000008a0000008a", 3771=>X"0000008a0000008a0000008a0000008a", 3772=>X"0000008a0000008a0000008a0000008a", 3773=>X"0000008a0000008a0000008a0000008a", 3774=>X"0000008a0000008a0000008a0000008a", 
3775=>X"0000008a0000008a0000008a0000008a", 3776=>X"00000089000000890000008a0000008a", 3777=>X"00000089000000890000008900000089", 3778=>X"00000089000000890000008900000089", 3779=>X"00000089000000890000008900000089", 
3780=>X"00000089000000890000008900000089", 3781=>X"00000089000000890000008900000089", 3782=>X"00000089000000890000008900000089", 3783=>X"00000089000000890000008900000089", 3784=>X"00000089000000890000008900000089", 
3785=>X"00000089000000890000008900000089", 3786=>X"00000089000000890000008900000089", 3787=>X"00000089000000890000008900000089", 3788=>X"00000089000000890000008900000089", 3789=>X"00000089000000890000008900000089", 
3790=>X"00000088000000880000008800000089", 3791=>X"00000088000000880000008800000088", 3792=>X"00000088000000880000008800000088", 3793=>X"00000088000000880000008800000088", 3794=>X"00000088000000880000008800000088", 
3795=>X"00000088000000880000008800000088", 3796=>X"00000088000000880000008800000088", 3797=>X"00000088000000880000008800000088", 3798=>X"00000088000000880000008800000088", 3799=>X"00000088000000880000008800000088", 
3800=>X"00000088000000880000008800000088", 3801=>X"00000088000000880000008800000088", 3802=>X"00000088000000880000008800000088", 3803=>X"00000088000000880000008800000088", 3804=>X"00000087000000870000008800000088", 
3805=>X"00000087000000870000008700000087", 3806=>X"00000087000000870000008700000087", 3807=>X"00000087000000870000008700000087", 3808=>X"00000087000000870000008700000087", 3809=>X"00000087000000870000008700000087", 
3810=>X"00000087000000870000008700000087", 3811=>X"00000087000000870000008700000087", 3812=>X"00000087000000870000008700000087", 3813=>X"00000087000000870000008700000087", 3814=>X"00000087000000870000008700000087", 
3815=>X"00000087000000870000008700000087", 3816=>X"00000087000000870000008700000087", 3817=>X"00000087000000870000008700000087", 3818=>X"00000087000000870000008700000087", 3819=>X"00000086000000860000008600000086", 
3820=>X"00000086000000860000008600000086", 3821=>X"00000086000000860000008600000086", 3822=>X"00000086000000860000008600000086", 3823=>X"00000086000000860000008600000086", 3824=>X"00000086000000860000008600000086", 
3825=>X"00000086000000860000008600000086", 3826=>X"00000086000000860000008600000086", 3827=>X"00000086000000860000008600000086", 3828=>X"00000086000000860000008600000086", 3829=>X"00000086000000860000008600000086", 
3830=>X"00000086000000860000008600000086", 3831=>X"00000086000000860000008600000086", 3832=>X"00000086000000860000008600000086", 3833=>X"00000085000000850000008600000086", 3834=>X"00000085000000850000008500000085", 
3835=>X"00000085000000850000008500000085", 3836=>X"00000085000000850000008500000085", 3837=>X"00000085000000850000008500000085", 3838=>X"00000085000000850000008500000085", 3839=>X"00000085000000850000008500000085", 
3840=>X"00000085000000850000008500000085", 3841=>X"00000085000000850000008500000085", 3842=>X"00000085000000850000008500000085", 3843=>X"00000085000000850000008500000085", 3844=>X"00000085000000850000008500000085", 
3845=>X"00000085000000850000008500000085", 3846=>X"00000085000000850000008500000085", 3847=>X"00000085000000850000008500000085", 3848=>X"00000084000000840000008400000085", 3849=>X"00000084000000840000008400000084", 
3850=>X"00000084000000840000008400000084", 3851=>X"00000084000000840000008400000084", 3852=>X"00000084000000840000008400000084", 3853=>X"00000084000000840000008400000084", 3854=>X"00000084000000840000008400000084", 
3855=>X"00000084000000840000008400000084", 3856=>X"00000084000000840000008400000084", 3857=>X"00000084000000840000008400000084", 3858=>X"00000084000000840000008400000084", 3859=>X"00000084000000840000008400000084", 
3860=>X"00000084000000840000008400000084", 3861=>X"00000084000000840000008400000084", 3862=>X"00000084000000840000008400000084", 3863=>X"00000083000000830000008300000084", 3864=>X"00000083000000830000008300000083", 
3865=>X"00000083000000830000008300000083", 3866=>X"00000083000000830000008300000083", 3867=>X"00000083000000830000008300000083", 3868=>X"00000083000000830000008300000083", 3869=>X"00000083000000830000008300000083", 
3870=>X"00000083000000830000008300000083", 3871=>X"00000083000000830000008300000083", 3872=>X"00000083000000830000008300000083", 3873=>X"00000083000000830000008300000083", 3874=>X"00000083000000830000008300000083", 
3875=>X"00000083000000830000008300000083", 3876=>X"00000083000000830000008300000083", 3877=>X"00000083000000830000008300000083", 3878=>X"00000082000000830000008300000083", 3879=>X"00000082000000820000008200000082", 
3880=>X"00000082000000820000008200000082", 3881=>X"00000082000000820000008200000082", 3882=>X"00000082000000820000008200000082", 3883=>X"00000082000000820000008200000082", 3884=>X"00000082000000820000008200000082", 
3885=>X"00000082000000820000008200000082", 3886=>X"00000082000000820000008200000082", 3887=>X"00000082000000820000008200000082", 3888=>X"00000082000000820000008200000082", 3889=>X"00000082000000820000008200000082", 
3890=>X"00000082000000820000008200000082", 3891=>X"00000082000000820000008200000082", 3892=>X"00000082000000820000008200000082", 3893=>X"00000082000000820000008200000082", 3894=>X"00000081000000810000008100000082", 
3895=>X"00000081000000810000008100000081", 3896=>X"00000081000000810000008100000081", 3897=>X"00000081000000810000008100000081", 3898=>X"00000081000000810000008100000081", 3899=>X"00000081000000810000008100000081", 
3900=>X"00000081000000810000008100000081", 3901=>X"00000081000000810000008100000081", 3902=>X"00000081000000810000008100000081", 3903=>X"00000081000000810000008100000081", 3904=>X"00000081000000810000008100000081", 
3905=>X"00000081000000810000008100000081", 3906=>X"00000081000000810000008100000081", 3907=>X"00000081000000810000008100000081", 3908=>X"00000081000000810000008100000081", 3909=>X"00000081000000810000008100000081", 
3910=>X"00000080000000800000008000000080", 3911=>X"00000080000000800000008000000080", 3912=>X"00000080000000800000008000000080", 3913=>X"00000080000000800000008000000080", 3914=>X"00000080000000800000008000000080", 
3915=>X"00000080000000800000008000000080", 3916=>X"00000080000000800000008000000080", 3917=>X"00000080000000800000008000000080", 3918=>X"00000080000000800000008000000080", 3919=>X"00000080000000800000008000000080", 
3920=>X"00000080000000800000008000000080", 3921=>X"00000080000000800000008000000080", 3922=>X"00000080000000800000008000000080", 3923=>X"00000080000000800000008000000080", 3924=>X"00000080000000800000008000000080", 
3925=>X"00000080000000800000008000000080", 3926=>X"0000007f0000007f0000007f0000007f", 3927=>X"0000007f0000007f0000007f0000007f", 3928=>X"0000007f0000007f0000007f0000007f", 3929=>X"0000007f0000007f0000007f0000007f", 
3930=>X"0000007f0000007f0000007f0000007f", 3931=>X"0000007f0000007f0000007f0000007f", 3932=>X"0000007f0000007f0000007f0000007f", 3933=>X"0000007f0000007f0000007f0000007f", 3934=>X"0000007f0000007f0000007f0000007f", 
3935=>X"0000007f0000007f0000007f0000007f", 3936=>X"0000007f0000007f0000007f0000007f", 3937=>X"0000007f0000007f0000007f0000007f", 3938=>X"0000007f0000007f0000007f0000007f", 3939=>X"0000007f0000007f0000007f0000007f", 
3940=>X"0000007f0000007f0000007f0000007f", 3941=>X"0000007f0000007f0000007f0000007f", 3942=>X"0000007e0000007e0000007e0000007f", 3943=>X"0000007e0000007e0000007e0000007e", 3944=>X"0000007e0000007e0000007e0000007e", 
3945=>X"0000007e0000007e0000007e0000007e", 3946=>X"0000007e0000007e0000007e0000007e", 3947=>X"0000007e0000007e0000007e0000007e", 3948=>X"0000007e0000007e0000007e0000007e", 3949=>X"0000007e0000007e0000007e0000007e", 
3950=>X"0000007e0000007e0000007e0000007e", 3951=>X"0000007e0000007e0000007e0000007e", 3952=>X"0000007e0000007e0000007e0000007e", 3953=>X"0000007e0000007e0000007e0000007e", 3954=>X"0000007e0000007e0000007e0000007e", 
3955=>X"0000007e0000007e0000007e0000007e", 3956=>X"0000007e0000007e0000007e0000007e", 3957=>X"0000007e0000007e0000007e0000007e", 3958=>X"0000007d0000007e0000007e0000007e", 3959=>X"0000007d0000007d0000007d0000007d", 
3960=>X"0000007d0000007d0000007d0000007d", 3961=>X"0000007d0000007d0000007d0000007d", 3962=>X"0000007d0000007d0000007d0000007d", 3963=>X"0000007d0000007d0000007d0000007d", 3964=>X"0000007d0000007d0000007d0000007d", 
3965=>X"0000007d0000007d0000007d0000007d", 3966=>X"0000007d0000007d0000007d0000007d", 3967=>X"0000007d0000007d0000007d0000007d", 3968=>X"0000007d0000007d0000007d0000007d", 3969=>X"0000007d0000007d0000007d0000007d", 
3970=>X"0000007d0000007d0000007d0000007d", 3971=>X"0000007d0000007d0000007d0000007d", 3972=>X"0000007d0000007d0000007d0000007d", 3973=>X"0000007d0000007d0000007d0000007d", 3974=>X"0000007d0000007d0000007d0000007d", 
3975=>X"0000007c0000007c0000007d0000007d", 3976=>X"0000007c0000007c0000007c0000007c", 3977=>X"0000007c0000007c0000007c0000007c", 3978=>X"0000007c0000007c0000007c0000007c", 3979=>X"0000007c0000007c0000007c0000007c", 
3980=>X"0000007c0000007c0000007c0000007c", 3981=>X"0000007c0000007c0000007c0000007c", 3982=>X"0000007c0000007c0000007c0000007c", 3983=>X"0000007c0000007c0000007c0000007c", 3984=>X"0000007c0000007c0000007c0000007c", 
3985=>X"0000007c0000007c0000007c0000007c", 3986=>X"0000007c0000007c0000007c0000007c", 3987=>X"0000007c0000007c0000007c0000007c", 3988=>X"0000007c0000007c0000007c0000007c", 3989=>X"0000007c0000007c0000007c0000007c", 
3990=>X"0000007c0000007c0000007c0000007c", 3991=>X"0000007c0000007c0000007c0000007c", 3992=>X"0000007b0000007b0000007c0000007c", 3993=>X"0000007b0000007b0000007b0000007b", 3994=>X"0000007b0000007b0000007b0000007b", 
3995=>X"0000007b0000007b0000007b0000007b", 3996=>X"0000007b0000007b0000007b0000007b", 3997=>X"0000007b0000007b0000007b0000007b", 3998=>X"0000007b0000007b0000007b0000007b", 3999=>X"0000007b0000007b0000007b0000007b", 
4000=>X"0000007b0000007b0000007b0000007b", 4001=>X"0000007b0000007b0000007b0000007b", 4002=>X"0000007b0000007b0000007b0000007b", 4003=>X"0000007b0000007b0000007b0000007b", 4004=>X"0000007b0000007b0000007b0000007b", 
4005=>X"0000007b0000007b0000007b0000007b", 4006=>X"0000007b0000007b0000007b0000007b", 4007=>X"0000007b0000007b0000007b0000007b", 4008=>X"0000007b0000007b0000007b0000007b", 4009=>X"0000007a0000007b0000007b0000007b", 
4010=>X"0000007a0000007a0000007a0000007a", 4011=>X"0000007a0000007a0000007a0000007a", 4012=>X"0000007a0000007a0000007a0000007a", 4013=>X"0000007a0000007a0000007a0000007a", 4014=>X"0000007a0000007a0000007a0000007a", 
4015=>X"0000007a0000007a0000007a0000007a", 4016=>X"0000007a0000007a0000007a0000007a", 4017=>X"0000007a0000007a0000007a0000007a", 4018=>X"0000007a0000007a0000007a0000007a", 4019=>X"0000007a0000007a0000007a0000007a", 
4020=>X"0000007a0000007a0000007a0000007a", 4021=>X"0000007a0000007a0000007a0000007a", 4022=>X"0000007a0000007a0000007a0000007a", 4023=>X"0000007a0000007a0000007a0000007a", 4024=>X"0000007a0000007a0000007a0000007a", 
4025=>X"0000007a0000007a0000007a0000007a", 4026=>X"0000007a0000007a0000007a0000007a", 4027=>X"00000079000000790000007a0000007a", 4028=>X"00000079000000790000007900000079", 4029=>X"00000079000000790000007900000079", 
4030=>X"00000079000000790000007900000079", 4031=>X"00000079000000790000007900000079", 4032=>X"00000079000000790000007900000079", 4033=>X"00000079000000790000007900000079", 4034=>X"00000079000000790000007900000079", 
4035=>X"00000079000000790000007900000079", 4036=>X"00000079000000790000007900000079", 4037=>X"00000079000000790000007900000079", 4038=>X"00000079000000790000007900000079", 4039=>X"00000079000000790000007900000079", 
4040=>X"00000079000000790000007900000079", 4041=>X"00000079000000790000007900000079", 4042=>X"00000079000000790000007900000079", 4043=>X"00000079000000790000007900000079", 4044=>X"00000079000000790000007900000079", 
4045=>X"00000078000000780000007800000079", 4046=>X"00000078000000780000007800000078", 4047=>X"00000078000000780000007800000078", 4048=>X"00000078000000780000007800000078", 4049=>X"00000078000000780000007800000078", 
4050=>X"00000078000000780000007800000078", 4051=>X"00000078000000780000007800000078", 4052=>X"00000078000000780000007800000078", 4053=>X"00000078000000780000007800000078", 4054=>X"00000078000000780000007800000078", 
4055=>X"00000078000000780000007800000078", 4056=>X"00000078000000780000007800000078", 4057=>X"00000078000000780000007800000078", 4058=>X"00000078000000780000007800000078", 4059=>X"00000078000000780000007800000078", 
4060=>X"00000078000000780000007800000078", 4061=>X"00000078000000780000007800000078", 4062=>X"00000078000000780000007800000078", 4063=>X"00000077000000770000007800000078", 4064=>X"00000077000000770000007700000077", 
4065=>X"00000077000000770000007700000077", 4066=>X"00000077000000770000007700000077", 4067=>X"00000077000000770000007700000077", 4068=>X"00000077000000770000007700000077", 4069=>X"00000077000000770000007700000077", 
4070=>X"00000077000000770000007700000077", 4071=>X"00000077000000770000007700000077", 4072=>X"00000077000000770000007700000077", 4073=>X"00000077000000770000007700000077", 4074=>X"00000077000000770000007700000077", 
4075=>X"00000077000000770000007700000077", 4076=>X"00000077000000770000007700000077", 4077=>X"00000077000000770000007700000077", 4078=>X"00000077000000770000007700000077", 4079=>X"00000077000000770000007700000077", 
4080=>X"00000077000000770000007700000077", 4081=>X"00000077000000770000007700000077", 4082=>X"00000076000000760000007600000076", 4083=>X"00000076000000760000007600000076", 4084=>X"00000076000000760000007600000076", 
4085=>X"00000076000000760000007600000076", 4086=>X"00000076000000760000007600000076", 4087=>X"00000076000000760000007600000076", 4088=>X"00000076000000760000007600000076", 4089=>X"00000076000000760000007600000076", 
4090=>X"00000076000000760000007600000076", 4091=>X"00000076000000760000007600000076", 4092=>X"00000076000000760000007600000076", 4093=>X"00000076000000760000007600000076", 4094=>X"00000076000000760000007600000076", 
4095=>X"00000076000000760000007600000076", 4096=>X"00000076000000760000007600000076", 4097=>X"00000076000000760000007600000076", 4098=>X"00000076000000760000007600000076", 4099=>X"00000076000000760000007600000076", 
4100=>X"00000076000000760000007600000076", 4101=>X"00000075000000750000007500000075", 4102=>X"00000075000000750000007500000075", 4103=>X"00000075000000750000007500000075", 4104=>X"00000075000000750000007500000075", 
4105=>X"00000075000000750000007500000075", 4106=>X"00000075000000750000007500000075", 4107=>X"00000075000000750000007500000075", 4108=>X"00000075000000750000007500000075", 4109=>X"00000075000000750000007500000075", 
4110=>X"00000075000000750000007500000075", 4111=>X"00000075000000750000007500000075", 4112=>X"00000075000000750000007500000075", 4113=>X"00000075000000750000007500000075", 4114=>X"00000075000000750000007500000075", 
4115=>X"00000075000000750000007500000075", 4116=>X"00000075000000750000007500000075", 4117=>X"00000075000000750000007500000075", 4118=>X"00000075000000750000007500000075", 4119=>X"00000075000000750000007500000075", 
4120=>X"00000074000000740000007400000074", 4121=>X"00000074000000740000007400000074", 4122=>X"00000074000000740000007400000074", 4123=>X"00000074000000740000007400000074", 4124=>X"00000074000000740000007400000074", 
4125=>X"00000074000000740000007400000074", 4126=>X"00000074000000740000007400000074", 4127=>X"00000074000000740000007400000074", 4128=>X"00000074000000740000007400000074", 4129=>X"00000074000000740000007400000074", 
4130=>X"00000074000000740000007400000074", 4131=>X"00000074000000740000007400000074", 4132=>X"00000074000000740000007400000074", 4133=>X"00000074000000740000007400000074", 4134=>X"00000074000000740000007400000074", 
4135=>X"00000074000000740000007400000074", 4136=>X"00000074000000740000007400000074", 4137=>X"00000074000000740000007400000074", 4138=>X"00000074000000740000007400000074", 4139=>X"00000073000000730000007400000074", 
4140=>X"00000073000000730000007300000073", 4141=>X"00000073000000730000007300000073", 4142=>X"00000073000000730000007300000073", 4143=>X"00000073000000730000007300000073", 4144=>X"00000073000000730000007300000073", 
4145=>X"00000073000000730000007300000073", 4146=>X"00000073000000730000007300000073", 4147=>X"00000073000000730000007300000073", 4148=>X"00000073000000730000007300000073", 4149=>X"00000073000000730000007300000073", 
4150=>X"00000073000000730000007300000073", 4151=>X"00000073000000730000007300000073", 4152=>X"00000073000000730000007300000073", 4153=>X"00000073000000730000007300000073", 4154=>X"00000073000000730000007300000073", 
4155=>X"00000073000000730000007300000073", 4156=>X"00000073000000730000007300000073", 4157=>X"00000073000000730000007300000073", 4158=>X"00000073000000730000007300000073", 4159=>X"00000072000000720000007200000073", 
4160=>X"00000072000000720000007200000072", 4161=>X"00000072000000720000007200000072", 4162=>X"00000072000000720000007200000072", 4163=>X"00000072000000720000007200000072", 4164=>X"00000072000000720000007200000072", 
4165=>X"00000072000000720000007200000072", 4166=>X"00000072000000720000007200000072", 4167=>X"00000072000000720000007200000072", 4168=>X"00000072000000720000007200000072", 4169=>X"00000072000000720000007200000072", 
4170=>X"00000072000000720000007200000072", 4171=>X"00000072000000720000007200000072", 4172=>X"00000072000000720000007200000072", 4173=>X"00000072000000720000007200000072", 4174=>X"00000072000000720000007200000072", 
4175=>X"00000072000000720000007200000072", 4176=>X"00000072000000720000007200000072", 4177=>X"00000072000000720000007200000072", 4178=>X"00000072000000720000007200000072", 4179=>X"00000071000000710000007200000072", 
4180=>X"00000071000000710000007100000071", 4181=>X"00000071000000710000007100000071", 4182=>X"00000071000000710000007100000071", 4183=>X"00000071000000710000007100000071", 4184=>X"00000071000000710000007100000071", 
4185=>X"00000071000000710000007100000071", 4186=>X"00000071000000710000007100000071", 4187=>X"00000071000000710000007100000071", 4188=>X"00000071000000710000007100000071", 4189=>X"00000071000000710000007100000071", 
4190=>X"00000071000000710000007100000071", 4191=>X"00000071000000710000007100000071", 4192=>X"00000071000000710000007100000071", 4193=>X"00000071000000710000007100000071", 4194=>X"00000071000000710000007100000071", 
4195=>X"00000071000000710000007100000071", 4196=>X"00000071000000710000007100000071", 4197=>X"00000071000000710000007100000071", 4198=>X"00000071000000710000007100000071", 4199=>X"00000071000000710000007100000071", 
4200=>X"00000070000000700000007000000070", 4201=>X"00000070000000700000007000000070", 4202=>X"00000070000000700000007000000070", 4203=>X"00000070000000700000007000000070", 4204=>X"00000070000000700000007000000070", 
4205=>X"00000070000000700000007000000070", 4206=>X"00000070000000700000007000000070", 4207=>X"00000070000000700000007000000070", 4208=>X"00000070000000700000007000000070", 4209=>X"00000070000000700000007000000070", 
4210=>X"00000070000000700000007000000070", 4211=>X"00000070000000700000007000000070", 4212=>X"00000070000000700000007000000070", 4213=>X"00000070000000700000007000000070", 4214=>X"00000070000000700000007000000070", 
4215=>X"00000070000000700000007000000070", 4216=>X"00000070000000700000007000000070", 4217=>X"00000070000000700000007000000070", 4218=>X"00000070000000700000007000000070", 4219=>X"00000070000000700000007000000070", 
4220=>X"00000070000000700000007000000070", 4221=>X"0000006f0000006f0000006f0000006f", 4222=>X"0000006f0000006f0000006f0000006f", 4223=>X"0000006f0000006f0000006f0000006f", 4224=>X"0000006f0000006f0000006f0000006f", 
4225=>X"0000006f0000006f0000006f0000006f", 4226=>X"0000006f0000006f0000006f0000006f", 4227=>X"0000006f0000006f0000006f0000006f", 4228=>X"0000006f0000006f0000006f0000006f", 4229=>X"0000006f0000006f0000006f0000006f", 
4230=>X"0000006f0000006f0000006f0000006f", 4231=>X"0000006f0000006f0000006f0000006f", 4232=>X"0000006f0000006f0000006f0000006f", 4233=>X"0000006f0000006f0000006f0000006f", 4234=>X"0000006f0000006f0000006f0000006f", 
4235=>X"0000006f0000006f0000006f0000006f", 4236=>X"0000006f0000006f0000006f0000006f", 4237=>X"0000006f0000006f0000006f0000006f", 4238=>X"0000006f0000006f0000006f0000006f", 4239=>X"0000006f0000006f0000006f0000006f", 
4240=>X"0000006f0000006f0000006f0000006f", 4241=>X"0000006f0000006f0000006f0000006f", 4242=>X"0000006e0000006e0000006e0000006f", 4243=>X"0000006e0000006e0000006e0000006e", 4244=>X"0000006e0000006e0000006e0000006e", 
4245=>X"0000006e0000006e0000006e0000006e", 4246=>X"0000006e0000006e0000006e0000006e", 4247=>X"0000006e0000006e0000006e0000006e", 4248=>X"0000006e0000006e0000006e0000006e", 4249=>X"0000006e0000006e0000006e0000006e", 
4250=>X"0000006e0000006e0000006e0000006e", 4251=>X"0000006e0000006e0000006e0000006e", 4252=>X"0000006e0000006e0000006e0000006e", 4253=>X"0000006e0000006e0000006e0000006e", 4254=>X"0000006e0000006e0000006e0000006e", 
4255=>X"0000006e0000006e0000006e0000006e", 4256=>X"0000006e0000006e0000006e0000006e", 4257=>X"0000006e0000006e0000006e0000006e", 4258=>X"0000006e0000006e0000006e0000006e", 4259=>X"0000006e0000006e0000006e0000006e", 
4260=>X"0000006e0000006e0000006e0000006e", 4261=>X"0000006e0000006e0000006e0000006e", 4262=>X"0000006e0000006e0000006e0000006e", 4263=>X"0000006e0000006e0000006e0000006e", 4264=>X"0000006d0000006d0000006d0000006d", 
4265=>X"0000006d0000006d0000006d0000006d", 4266=>X"0000006d0000006d0000006d0000006d", 4267=>X"0000006d0000006d0000006d0000006d", 4268=>X"0000006d0000006d0000006d0000006d", 4269=>X"0000006d0000006d0000006d0000006d", 
4270=>X"0000006d0000006d0000006d0000006d", 4271=>X"0000006d0000006d0000006d0000006d", 4272=>X"0000006d0000006d0000006d0000006d", 4273=>X"0000006d0000006d0000006d0000006d", 4274=>X"0000006d0000006d0000006d0000006d", 
4275=>X"0000006d0000006d0000006d0000006d", 4276=>X"0000006d0000006d0000006d0000006d", 4277=>X"0000006d0000006d0000006d0000006d", 4278=>X"0000006d0000006d0000006d0000006d", 4279=>X"0000006d0000006d0000006d0000006d", 
4280=>X"0000006d0000006d0000006d0000006d", 4281=>X"0000006d0000006d0000006d0000006d", 4282=>X"0000006d0000006d0000006d0000006d", 4283=>X"0000006d0000006d0000006d0000006d", 4284=>X"0000006d0000006d0000006d0000006d", 
4285=>X"0000006d0000006d0000006d0000006d", 4286=>X"0000006c0000006c0000006c0000006c", 4287=>X"0000006c0000006c0000006c0000006c", 4288=>X"0000006c0000006c0000006c0000006c", 4289=>X"0000006c0000006c0000006c0000006c", 
4290=>X"0000006c0000006c0000006c0000006c", 4291=>X"0000006c0000006c0000006c0000006c", 4292=>X"0000006c0000006c0000006c0000006c", 4293=>X"0000006c0000006c0000006c0000006c", 4294=>X"0000006c0000006c0000006c0000006c", 
4295=>X"0000006c0000006c0000006c0000006c", 4296=>X"0000006c0000006c0000006c0000006c", 4297=>X"0000006c0000006c0000006c0000006c", 4298=>X"0000006c0000006c0000006c0000006c", 4299=>X"0000006c0000006c0000006c0000006c", 
4300=>X"0000006c0000006c0000006c0000006c", 4301=>X"0000006c0000006c0000006c0000006c", 4302=>X"0000006c0000006c0000006c0000006c", 4303=>X"0000006c0000006c0000006c0000006c", 4304=>X"0000006c0000006c0000006c0000006c", 
4305=>X"0000006c0000006c0000006c0000006c", 4306=>X"0000006c0000006c0000006c0000006c", 4307=>X"0000006c0000006c0000006c0000006c", 4308=>X"0000006b0000006b0000006c0000006c", 4309=>X"0000006b0000006b0000006b0000006b", 
4310=>X"0000006b0000006b0000006b0000006b", 4311=>X"0000006b0000006b0000006b0000006b", 4312=>X"0000006b0000006b0000006b0000006b", 4313=>X"0000006b0000006b0000006b0000006b", 4314=>X"0000006b0000006b0000006b0000006b", 
4315=>X"0000006b0000006b0000006b0000006b", 4316=>X"0000006b0000006b0000006b0000006b", 4317=>X"0000006b0000006b0000006b0000006b", 4318=>X"0000006b0000006b0000006b0000006b", 4319=>X"0000006b0000006b0000006b0000006b", 
4320=>X"0000006b0000006b0000006b0000006b", 4321=>X"0000006b0000006b0000006b0000006b", 4322=>X"0000006b0000006b0000006b0000006b", 4323=>X"0000006b0000006b0000006b0000006b", 4324=>X"0000006b0000006b0000006b0000006b", 
4325=>X"0000006b0000006b0000006b0000006b", 4326=>X"0000006b0000006b0000006b0000006b", 4327=>X"0000006b0000006b0000006b0000006b", 4328=>X"0000006b0000006b0000006b0000006b", 4329=>X"0000006b0000006b0000006b0000006b", 
4330=>X"0000006b0000006b0000006b0000006b", 4331=>X"0000006a0000006a0000006a0000006b", 4332=>X"0000006a0000006a0000006a0000006a", 4333=>X"0000006a0000006a0000006a0000006a", 4334=>X"0000006a0000006a0000006a0000006a", 
4335=>X"0000006a0000006a0000006a0000006a", 4336=>X"0000006a0000006a0000006a0000006a", 4337=>X"0000006a0000006a0000006a0000006a", 4338=>X"0000006a0000006a0000006a0000006a", 4339=>X"0000006a0000006a0000006a0000006a", 
4340=>X"0000006a0000006a0000006a0000006a", 4341=>X"0000006a0000006a0000006a0000006a", 4342=>X"0000006a0000006a0000006a0000006a", 4343=>X"0000006a0000006a0000006a0000006a", 4344=>X"0000006a0000006a0000006a0000006a", 
4345=>X"0000006a0000006a0000006a0000006a", 4346=>X"0000006a0000006a0000006a0000006a", 4347=>X"0000006a0000006a0000006a0000006a", 4348=>X"0000006a0000006a0000006a0000006a", 4349=>X"0000006a0000006a0000006a0000006a", 
4350=>X"0000006a0000006a0000006a0000006a", 4351=>X"0000006a0000006a0000006a0000006a", 4352=>X"0000006a0000006a0000006a0000006a", 4353=>X"0000006a0000006a0000006a0000006a", 4354=>X"000000690000006a0000006a0000006a", 
4355=>X"00000069000000690000006900000069", 4356=>X"00000069000000690000006900000069", 4357=>X"00000069000000690000006900000069", 4358=>X"00000069000000690000006900000069", 4359=>X"00000069000000690000006900000069", 
4360=>X"00000069000000690000006900000069", 4361=>X"00000069000000690000006900000069", 4362=>X"00000069000000690000006900000069", 4363=>X"00000069000000690000006900000069", 4364=>X"00000069000000690000006900000069", 
4365=>X"00000069000000690000006900000069", 4366=>X"00000069000000690000006900000069", 4367=>X"00000069000000690000006900000069", 4368=>X"00000069000000690000006900000069", 4369=>X"00000069000000690000006900000069", 
4370=>X"00000069000000690000006900000069", 4371=>X"00000069000000690000006900000069", 4372=>X"00000069000000690000006900000069", 4373=>X"00000069000000690000006900000069", 4374=>X"00000069000000690000006900000069", 
4375=>X"00000069000000690000006900000069", 4376=>X"00000069000000690000006900000069", 4377=>X"00000069000000690000006900000069", 4378=>X"00000068000000680000006900000069", 4379=>X"00000068000000680000006800000068", 
4380=>X"00000068000000680000006800000068", 4381=>X"00000068000000680000006800000068", 4382=>X"00000068000000680000006800000068", 4383=>X"00000068000000680000006800000068", 4384=>X"00000068000000680000006800000068", 
4385=>X"00000068000000680000006800000068", 4386=>X"00000068000000680000006800000068", 4387=>X"00000068000000680000006800000068", 4388=>X"00000068000000680000006800000068", 4389=>X"00000068000000680000006800000068", 
4390=>X"00000068000000680000006800000068", 4391=>X"00000068000000680000006800000068", 4392=>X"00000068000000680000006800000068", 4393=>X"00000068000000680000006800000068", 4394=>X"00000068000000680000006800000068", 
4395=>X"00000068000000680000006800000068", 4396=>X"00000068000000680000006800000068", 4397=>X"00000068000000680000006800000068", 4398=>X"00000068000000680000006800000068", 4399=>X"00000068000000680000006800000068", 
4400=>X"00000068000000680000006800000068", 4401=>X"00000068000000680000006800000068", 4402=>X"00000067000000680000006800000068", 4403=>X"00000067000000670000006700000067", 4404=>X"00000067000000670000006700000067", 
4405=>X"00000067000000670000006700000067", 4406=>X"00000067000000670000006700000067", 4407=>X"00000067000000670000006700000067", 4408=>X"00000067000000670000006700000067", 4409=>X"00000067000000670000006700000067", 
4410=>X"00000067000000670000006700000067", 4411=>X"00000067000000670000006700000067", 4412=>X"00000067000000670000006700000067", 4413=>X"00000067000000670000006700000067", 4414=>X"00000067000000670000006700000067", 
4415=>X"00000067000000670000006700000067", 4416=>X"00000067000000670000006700000067", 4417=>X"00000067000000670000006700000067", 4418=>X"00000067000000670000006700000067", 4419=>X"00000067000000670000006700000067", 
4420=>X"00000067000000670000006700000067", 4421=>X"00000067000000670000006700000067", 4422=>X"00000067000000670000006700000067", 4423=>X"00000067000000670000006700000067", 4424=>X"00000067000000670000006700000067", 
4425=>X"00000067000000670000006700000067", 4426=>X"00000067000000670000006700000067", 4427=>X"00000066000000660000006700000067", 4428=>X"00000066000000660000006600000066", 4429=>X"00000066000000660000006600000066", 
4430=>X"00000066000000660000006600000066", 4431=>X"00000066000000660000006600000066", 4432=>X"00000066000000660000006600000066", 4433=>X"00000066000000660000006600000066", 4434=>X"00000066000000660000006600000066", 
4435=>X"00000066000000660000006600000066", 4436=>X"00000066000000660000006600000066", 4437=>X"00000066000000660000006600000066", 4438=>X"00000066000000660000006600000066", 4439=>X"00000066000000660000006600000066", 
4440=>X"00000066000000660000006600000066", 4441=>X"00000066000000660000006600000066", 4442=>X"00000066000000660000006600000066", 4443=>X"00000066000000660000006600000066", 4444=>X"00000066000000660000006600000066", 
4445=>X"00000066000000660000006600000066", 4446=>X"00000066000000660000006600000066", 4447=>X"00000066000000660000006600000066", 4448=>X"00000066000000660000006600000066", 4449=>X"00000066000000660000006600000066", 
4450=>X"00000066000000660000006600000066", 4451=>X"00000066000000660000006600000066", 4452=>X"00000065000000650000006600000066", 4453=>X"00000065000000650000006500000065", 4454=>X"00000065000000650000006500000065", 
4455=>X"00000065000000650000006500000065", 4456=>X"00000065000000650000006500000065", 4457=>X"00000065000000650000006500000065", 4458=>X"00000065000000650000006500000065", 4459=>X"00000065000000650000006500000065", 
4460=>X"00000065000000650000006500000065", 4461=>X"00000065000000650000006500000065", 4462=>X"00000065000000650000006500000065", 4463=>X"00000065000000650000006500000065", 4464=>X"00000065000000650000006500000065", 
4465=>X"00000065000000650000006500000065", 4466=>X"00000065000000650000006500000065", 4467=>X"00000065000000650000006500000065", 4468=>X"00000065000000650000006500000065", 4469=>X"00000065000000650000006500000065", 
4470=>X"00000065000000650000006500000065", 4471=>X"00000065000000650000006500000065", 4472=>X"00000065000000650000006500000065", 4473=>X"00000065000000650000006500000065", 4474=>X"00000065000000650000006500000065", 
4475=>X"00000065000000650000006500000065", 4476=>X"00000065000000650000006500000065", 4477=>X"00000065000000650000006500000065", 4478=>X"00000064000000640000006400000065", 4479=>X"00000064000000640000006400000064", 
4480=>X"00000064000000640000006400000064", 4481=>X"00000064000000640000006400000064", 4482=>X"00000064000000640000006400000064", 4483=>X"00000064000000640000006400000064", 4484=>X"00000064000000640000006400000064", 
4485=>X"00000064000000640000006400000064", 4486=>X"00000064000000640000006400000064", 4487=>X"00000064000000640000006400000064", 4488=>X"00000064000000640000006400000064", 4489=>X"00000064000000640000006400000064", 
4490=>X"00000064000000640000006400000064", 4491=>X"00000064000000640000006400000064", 4492=>X"00000064000000640000006400000064", 4493=>X"00000064000000640000006400000064", 4494=>X"00000064000000640000006400000064", 
4495=>X"00000064000000640000006400000064", 4496=>X"00000064000000640000006400000064", 4497=>X"00000064000000640000006400000064", 4498=>X"00000064000000640000006400000064", 4499=>X"00000064000000640000006400000064", 
4500=>X"00000064000000640000006400000064", 4501=>X"00000064000000640000006400000064", 4502=>X"00000064000000640000006400000064", 4503=>X"00000064000000640000006400000064", 4504=>X"00000063000000630000006400000064", 
4505=>X"00000063000000630000006300000063", 4506=>X"00000063000000630000006300000063", 4507=>X"00000063000000630000006300000063", 4508=>X"00000063000000630000006300000063", 4509=>X"00000063000000630000006300000063", 
4510=>X"00000063000000630000006300000063", 4511=>X"00000063000000630000006300000063", 4512=>X"00000063000000630000006300000063", 4513=>X"00000063000000630000006300000063", 4514=>X"00000063000000630000006300000063", 
4515=>X"00000063000000630000006300000063", 4516=>X"00000063000000630000006300000063", 4517=>X"00000063000000630000006300000063", 4518=>X"00000063000000630000006300000063", 4519=>X"00000063000000630000006300000063", 
4520=>X"00000063000000630000006300000063", 4521=>X"00000063000000630000006300000063", 4522=>X"00000063000000630000006300000063", 4523=>X"00000063000000630000006300000063", 4524=>X"00000063000000630000006300000063", 
4525=>X"00000063000000630000006300000063", 4526=>X"00000063000000630000006300000063", 4527=>X"00000063000000630000006300000063", 4528=>X"00000063000000630000006300000063", 4529=>X"00000063000000630000006300000063", 
4530=>X"00000063000000630000006300000063", 4531=>X"00000062000000620000006200000063", 4532=>X"00000062000000620000006200000062", 4533=>X"00000062000000620000006200000062", 4534=>X"00000062000000620000006200000062", 
4535=>X"00000062000000620000006200000062", 4536=>X"00000062000000620000006200000062", 4537=>X"00000062000000620000006200000062", 4538=>X"00000062000000620000006200000062", 4539=>X"00000062000000620000006200000062", 
4540=>X"00000062000000620000006200000062", 4541=>X"00000062000000620000006200000062", 4542=>X"00000062000000620000006200000062", 4543=>X"00000062000000620000006200000062", 4544=>X"00000062000000620000006200000062", 
4545=>X"00000062000000620000006200000062", 4546=>X"00000062000000620000006200000062", 4547=>X"00000062000000620000006200000062", 4548=>X"00000062000000620000006200000062", 4549=>X"00000062000000620000006200000062", 
4550=>X"00000062000000620000006200000062", 4551=>X"00000062000000620000006200000062", 4552=>X"00000062000000620000006200000062", 4553=>X"00000062000000620000006200000062", 4554=>X"00000062000000620000006200000062", 
4555=>X"00000062000000620000006200000062", 4556=>X"00000062000000620000006200000062", 4557=>X"00000062000000620000006200000062", 4558=>X"00000061000000610000006200000062", 4559=>X"00000061000000610000006100000061", 
4560=>X"00000061000000610000006100000061", 4561=>X"00000061000000610000006100000061", 4562=>X"00000061000000610000006100000061", 4563=>X"00000061000000610000006100000061", 4564=>X"00000061000000610000006100000061", 
4565=>X"00000061000000610000006100000061", 4566=>X"00000061000000610000006100000061", 4567=>X"00000061000000610000006100000061", 4568=>X"00000061000000610000006100000061", 4569=>X"00000061000000610000006100000061", 
4570=>X"00000061000000610000006100000061", 4571=>X"00000061000000610000006100000061", 4572=>X"00000061000000610000006100000061", 4573=>X"00000061000000610000006100000061", 4574=>X"00000061000000610000006100000061", 
4575=>X"00000061000000610000006100000061", 4576=>X"00000061000000610000006100000061", 4577=>X"00000061000000610000006100000061", 4578=>X"00000061000000610000006100000061", 4579=>X"00000061000000610000006100000061", 
4580=>X"00000061000000610000006100000061", 4581=>X"00000061000000610000006100000061", 4582=>X"00000061000000610000006100000061", 4583=>X"00000061000000610000006100000061", 4584=>X"00000061000000610000006100000061", 
4585=>X"00000061000000610000006100000061", 4586=>X"00000060000000600000006100000061", 4587=>X"00000060000000600000006000000060", 4588=>X"00000060000000600000006000000060", 4589=>X"00000060000000600000006000000060", 
4590=>X"00000060000000600000006000000060", 4591=>X"00000060000000600000006000000060", 4592=>X"00000060000000600000006000000060", 4593=>X"00000060000000600000006000000060", 4594=>X"00000060000000600000006000000060", 
4595=>X"00000060000000600000006000000060", 4596=>X"00000060000000600000006000000060", 4597=>X"00000060000000600000006000000060", 4598=>X"00000060000000600000006000000060", 4599=>X"00000060000000600000006000000060", 
4600=>X"00000060000000600000006000000060", 4601=>X"00000060000000600000006000000060", 4602=>X"00000060000000600000006000000060", 4603=>X"00000060000000600000006000000060", 4604=>X"00000060000000600000006000000060", 
4605=>X"00000060000000600000006000000060", 4606=>X"00000060000000600000006000000060", 4607=>X"00000060000000600000006000000060", 4608=>X"00000060000000600000006000000060", 4609=>X"00000060000000600000006000000060", 
4610=>X"00000060000000600000006000000060", 4611=>X"00000060000000600000006000000060", 4612=>X"00000060000000600000006000000060", 4613=>X"00000060000000600000006000000060", 4614=>X"0000005f000000600000006000000060", 
4615=>X"0000005f0000005f0000005f0000005f", 4616=>X"0000005f0000005f0000005f0000005f", 4617=>X"0000005f0000005f0000005f0000005f", 4618=>X"0000005f0000005f0000005f0000005f", 4619=>X"0000005f0000005f0000005f0000005f", 
4620=>X"0000005f0000005f0000005f0000005f", 4621=>X"0000005f0000005f0000005f0000005f", 4622=>X"0000005f0000005f0000005f0000005f", 4623=>X"0000005f0000005f0000005f0000005f", 4624=>X"0000005f0000005f0000005f0000005f", 
4625=>X"0000005f0000005f0000005f0000005f", 4626=>X"0000005f0000005f0000005f0000005f", 4627=>X"0000005f0000005f0000005f0000005f", 4628=>X"0000005f0000005f0000005f0000005f", 4629=>X"0000005f0000005f0000005f0000005f", 
4630=>X"0000005f0000005f0000005f0000005f", 4631=>X"0000005f0000005f0000005f0000005f", 4632=>X"0000005f0000005f0000005f0000005f", 4633=>X"0000005f0000005f0000005f0000005f", 4634=>X"0000005f0000005f0000005f0000005f", 
4635=>X"0000005f0000005f0000005f0000005f", 4636=>X"0000005f0000005f0000005f0000005f", 4637=>X"0000005f0000005f0000005f0000005f", 4638=>X"0000005f0000005f0000005f0000005f", 4639=>X"0000005f0000005f0000005f0000005f", 
4640=>X"0000005f0000005f0000005f0000005f", 4641=>X"0000005f0000005f0000005f0000005f", 4642=>X"0000005f0000005f0000005f0000005f", 4643=>X"0000005f0000005f0000005f0000005f", 4644=>X"0000005e0000005e0000005e0000005e", 
4645=>X"0000005e0000005e0000005e0000005e", 4646=>X"0000005e0000005e0000005e0000005e", 4647=>X"0000005e0000005e0000005e0000005e", 4648=>X"0000005e0000005e0000005e0000005e", 4649=>X"0000005e0000005e0000005e0000005e", 
4650=>X"0000005e0000005e0000005e0000005e", 4651=>X"0000005e0000005e0000005e0000005e", 4652=>X"0000005e0000005e0000005e0000005e", 4653=>X"0000005e0000005e0000005e0000005e", 4654=>X"0000005e0000005e0000005e0000005e", 
4655=>X"0000005e0000005e0000005e0000005e", 4656=>X"0000005e0000005e0000005e0000005e", 4657=>X"0000005e0000005e0000005e0000005e", 4658=>X"0000005e0000005e0000005e0000005e", 4659=>X"0000005e0000005e0000005e0000005e", 
4660=>X"0000005e0000005e0000005e0000005e", 4661=>X"0000005e0000005e0000005e0000005e", 4662=>X"0000005e0000005e0000005e0000005e", 4663=>X"0000005e0000005e0000005e0000005e", 4664=>X"0000005e0000005e0000005e0000005e", 
4665=>X"0000005e0000005e0000005e0000005e", 4666=>X"0000005e0000005e0000005e0000005e", 4667=>X"0000005e0000005e0000005e0000005e", 4668=>X"0000005e0000005e0000005e0000005e", 4669=>X"0000005e0000005e0000005e0000005e", 
4670=>X"0000005e0000005e0000005e0000005e", 4671=>X"0000005e0000005e0000005e0000005e", 4672=>X"0000005e0000005e0000005e0000005e", 4673=>X"0000005d0000005d0000005e0000005e", 4674=>X"0000005d0000005d0000005d0000005d", 
4675=>X"0000005d0000005d0000005d0000005d", 4676=>X"0000005d0000005d0000005d0000005d", 4677=>X"0000005d0000005d0000005d0000005d", 4678=>X"0000005d0000005d0000005d0000005d", 4679=>X"0000005d0000005d0000005d0000005d", 
4680=>X"0000005d0000005d0000005d0000005d", 4681=>X"0000005d0000005d0000005d0000005d", 4682=>X"0000005d0000005d0000005d0000005d", 4683=>X"0000005d0000005d0000005d0000005d", 4684=>X"0000005d0000005d0000005d0000005d", 
4685=>X"0000005d0000005d0000005d0000005d", 4686=>X"0000005d0000005d0000005d0000005d", 4687=>X"0000005d0000005d0000005d0000005d", 4688=>X"0000005d0000005d0000005d0000005d", 4689=>X"0000005d0000005d0000005d0000005d", 
4690=>X"0000005d0000005d0000005d0000005d", 4691=>X"0000005d0000005d0000005d0000005d", 4692=>X"0000005d0000005d0000005d0000005d", 4693=>X"0000005d0000005d0000005d0000005d", 4694=>X"0000005d0000005d0000005d0000005d", 
4695=>X"0000005d0000005d0000005d0000005d", 4696=>X"0000005d0000005d0000005d0000005d", 4697=>X"0000005d0000005d0000005d0000005d", 4698=>X"0000005d0000005d0000005d0000005d", 4699=>X"0000005d0000005d0000005d0000005d", 
4700=>X"0000005d0000005d0000005d0000005d", 4701=>X"0000005d0000005d0000005d0000005d", 4702=>X"0000005d0000005d0000005d0000005d", 4703=>X"0000005c0000005d0000005d0000005d", 4704=>X"0000005c0000005c0000005c0000005c", 
4705=>X"0000005c0000005c0000005c0000005c", 4706=>X"0000005c0000005c0000005c0000005c", 4707=>X"0000005c0000005c0000005c0000005c", 4708=>X"0000005c0000005c0000005c0000005c", 4709=>X"0000005c0000005c0000005c0000005c", 
4710=>X"0000005c0000005c0000005c0000005c", 4711=>X"0000005c0000005c0000005c0000005c", 4712=>X"0000005c0000005c0000005c0000005c", 4713=>X"0000005c0000005c0000005c0000005c", 4714=>X"0000005c0000005c0000005c0000005c", 
4715=>X"0000005c0000005c0000005c0000005c", 4716=>X"0000005c0000005c0000005c0000005c", 4717=>X"0000005c0000005c0000005c0000005c", 4718=>X"0000005c0000005c0000005c0000005c", 4719=>X"0000005c0000005c0000005c0000005c", 
4720=>X"0000005c0000005c0000005c0000005c", 4721=>X"0000005c0000005c0000005c0000005c", 4722=>X"0000005c0000005c0000005c0000005c", 4723=>X"0000005c0000005c0000005c0000005c", 4724=>X"0000005c0000005c0000005c0000005c", 
4725=>X"0000005c0000005c0000005c0000005c", 4726=>X"0000005c0000005c0000005c0000005c", 4727=>X"0000005c0000005c0000005c0000005c", 4728=>X"0000005c0000005c0000005c0000005c", 4729=>X"0000005c0000005c0000005c0000005c", 
4730=>X"0000005c0000005c0000005c0000005c", 4731=>X"0000005c0000005c0000005c0000005c", 4732=>X"0000005c0000005c0000005c0000005c", 4733=>X"0000005c0000005c0000005c0000005c", 4734=>X"0000005b0000005c0000005c0000005c", 
4735=>X"0000005b0000005b0000005b0000005b", 4736=>X"0000005b0000005b0000005b0000005b", 4737=>X"0000005b0000005b0000005b0000005b", 4738=>X"0000005b0000005b0000005b0000005b", 4739=>X"0000005b0000005b0000005b0000005b", 
4740=>X"0000005b0000005b0000005b0000005b", 4741=>X"0000005b0000005b0000005b0000005b", 4742=>X"0000005b0000005b0000005b0000005b", 4743=>X"0000005b0000005b0000005b0000005b", 4744=>X"0000005b0000005b0000005b0000005b", 
4745=>X"0000005b0000005b0000005b0000005b", 4746=>X"0000005b0000005b0000005b0000005b", 4747=>X"0000005b0000005b0000005b0000005b", 4748=>X"0000005b0000005b0000005b0000005b", 4749=>X"0000005b0000005b0000005b0000005b", 
4750=>X"0000005b0000005b0000005b0000005b", 4751=>X"0000005b0000005b0000005b0000005b", 4752=>X"0000005b0000005b0000005b0000005b", 4753=>X"0000005b0000005b0000005b0000005b", 4754=>X"0000005b0000005b0000005b0000005b", 
4755=>X"0000005b0000005b0000005b0000005b", 4756=>X"0000005b0000005b0000005b0000005b", 4757=>X"0000005b0000005b0000005b0000005b", 4758=>X"0000005b0000005b0000005b0000005b", 4759=>X"0000005b0000005b0000005b0000005b", 
4760=>X"0000005b0000005b0000005b0000005b", 4761=>X"0000005b0000005b0000005b0000005b", 4762=>X"0000005b0000005b0000005b0000005b", 4763=>X"0000005b0000005b0000005b0000005b", 4764=>X"0000005b0000005b0000005b0000005b", 
4765=>X"0000005b0000005b0000005b0000005b", 4766=>X"0000005a0000005a0000005b0000005b", 4767=>X"0000005a0000005a0000005a0000005a", 4768=>X"0000005a0000005a0000005a0000005a", 4769=>X"0000005a0000005a0000005a0000005a", 
4770=>X"0000005a0000005a0000005a0000005a", 4771=>X"0000005a0000005a0000005a0000005a", 4772=>X"0000005a0000005a0000005a0000005a", 4773=>X"0000005a0000005a0000005a0000005a", 4774=>X"0000005a0000005a0000005a0000005a", 
4775=>X"0000005a0000005a0000005a0000005a", 4776=>X"0000005a0000005a0000005a0000005a", 4777=>X"0000005a0000005a0000005a0000005a", 4778=>X"0000005a0000005a0000005a0000005a", 4779=>X"0000005a0000005a0000005a0000005a", 
4780=>X"0000005a0000005a0000005a0000005a", 4781=>X"0000005a0000005a0000005a0000005a", 4782=>X"0000005a0000005a0000005a0000005a", 4783=>X"0000005a0000005a0000005a0000005a", 4784=>X"0000005a0000005a0000005a0000005a", 
4785=>X"0000005a0000005a0000005a0000005a", 4786=>X"0000005a0000005a0000005a0000005a", 4787=>X"0000005a0000005a0000005a0000005a", 4788=>X"0000005a0000005a0000005a0000005a", 4789=>X"0000005a0000005a0000005a0000005a", 
4790=>X"0000005a0000005a0000005a0000005a", 4791=>X"0000005a0000005a0000005a0000005a", 4792=>X"0000005a0000005a0000005a0000005a", 4793=>X"0000005a0000005a0000005a0000005a", 4794=>X"0000005a0000005a0000005a0000005a", 
4795=>X"0000005a0000005a0000005a0000005a", 4796=>X"0000005a0000005a0000005a0000005a", 4797=>X"0000005a0000005a0000005a0000005a", 4798=>X"000000590000005a0000005a0000005a", 4799=>X"00000059000000590000005900000059", 
4800=>X"00000059000000590000005900000059", 4801=>X"00000059000000590000005900000059", 4802=>X"00000059000000590000005900000059", 4803=>X"00000059000000590000005900000059", 4804=>X"00000059000000590000005900000059", 
4805=>X"00000059000000590000005900000059", 4806=>X"00000059000000590000005900000059", 4807=>X"00000059000000590000005900000059", 4808=>X"00000059000000590000005900000059", 4809=>X"00000059000000590000005900000059", 
4810=>X"00000059000000590000005900000059", 4811=>X"00000059000000590000005900000059", 4812=>X"00000059000000590000005900000059", 4813=>X"00000059000000590000005900000059", 4814=>X"00000059000000590000005900000059", 
4815=>X"00000059000000590000005900000059", 4816=>X"00000059000000590000005900000059", 4817=>X"00000059000000590000005900000059", 4818=>X"00000059000000590000005900000059", 4819=>X"00000059000000590000005900000059", 
4820=>X"00000059000000590000005900000059", 4821=>X"00000059000000590000005900000059", 4822=>X"00000059000000590000005900000059", 4823=>X"00000059000000590000005900000059", 4824=>X"00000059000000590000005900000059", 
4825=>X"00000059000000590000005900000059", 4826=>X"00000059000000590000005900000059", 4827=>X"00000059000000590000005900000059", 4828=>X"00000059000000590000005900000059", 4829=>X"00000059000000590000005900000059", 
4830=>X"00000059000000590000005900000059", 4831=>X"00000059000000590000005900000059", 4832=>X"00000058000000580000005800000058", 4833=>X"00000058000000580000005800000058", 4834=>X"00000058000000580000005800000058", 
4835=>X"00000058000000580000005800000058", 4836=>X"00000058000000580000005800000058", 4837=>X"00000058000000580000005800000058", 4838=>X"00000058000000580000005800000058", 4839=>X"00000058000000580000005800000058", 
4840=>X"00000058000000580000005800000058", 4841=>X"00000058000000580000005800000058", 4842=>X"00000058000000580000005800000058", 4843=>X"00000058000000580000005800000058", 4844=>X"00000058000000580000005800000058", 
4845=>X"00000058000000580000005800000058", 4846=>X"00000058000000580000005800000058", 4847=>X"00000058000000580000005800000058", 4848=>X"00000058000000580000005800000058", 4849=>X"00000058000000580000005800000058", 
4850=>X"00000058000000580000005800000058", 4851=>X"00000058000000580000005800000058", 4852=>X"00000058000000580000005800000058", 4853=>X"00000058000000580000005800000058", 4854=>X"00000058000000580000005800000058", 
4855=>X"00000058000000580000005800000058", 4856=>X"00000058000000580000005800000058", 4857=>X"00000058000000580000005800000058", 4858=>X"00000058000000580000005800000058", 4859=>X"00000058000000580000005800000058", 
4860=>X"00000058000000580000005800000058", 4861=>X"00000058000000580000005800000058", 4862=>X"00000058000000580000005800000058", 4863=>X"00000058000000580000005800000058", 4864=>X"00000058000000580000005800000058", 
4865=>X"00000057000000580000005800000058", 4866=>X"00000057000000570000005700000057", 4867=>X"00000057000000570000005700000057", 4868=>X"00000057000000570000005700000057", 4869=>X"00000057000000570000005700000057", 
4870=>X"00000057000000570000005700000057", 4871=>X"00000057000000570000005700000057", 4872=>X"00000057000000570000005700000057", 4873=>X"00000057000000570000005700000057", 4874=>X"00000057000000570000005700000057", 
4875=>X"00000057000000570000005700000057", 4876=>X"00000057000000570000005700000057", 4877=>X"00000057000000570000005700000057", 4878=>X"00000057000000570000005700000057", 4879=>X"00000057000000570000005700000057", 
4880=>X"00000057000000570000005700000057", 4881=>X"00000057000000570000005700000057", 4882=>X"00000057000000570000005700000057", 4883=>X"00000057000000570000005700000057", 4884=>X"00000057000000570000005700000057", 
4885=>X"00000057000000570000005700000057", 4886=>X"00000057000000570000005700000057", 4887=>X"00000057000000570000005700000057", 4888=>X"00000057000000570000005700000057", 4889=>X"00000057000000570000005700000057", 
4890=>X"00000057000000570000005700000057", 4891=>X"00000057000000570000005700000057", 4892=>X"00000057000000570000005700000057", 4893=>X"00000057000000570000005700000057", 4894=>X"00000057000000570000005700000057", 
4895=>X"00000057000000570000005700000057", 4896=>X"00000057000000570000005700000057", 4897=>X"00000057000000570000005700000057", 4898=>X"00000057000000570000005700000057", 4899=>X"00000057000000570000005700000057", 
4900=>X"00000056000000560000005700000057", 4901=>X"00000056000000560000005600000056", 4902=>X"00000056000000560000005600000056", 4903=>X"00000056000000560000005600000056", 4904=>X"00000056000000560000005600000056", 
4905=>X"00000056000000560000005600000056", 4906=>X"00000056000000560000005600000056", 4907=>X"00000056000000560000005600000056", 4908=>X"00000056000000560000005600000056", 4909=>X"00000056000000560000005600000056", 
4910=>X"00000056000000560000005600000056", 4911=>X"00000056000000560000005600000056", 4912=>X"00000056000000560000005600000056", 4913=>X"00000056000000560000005600000056", 4914=>X"00000056000000560000005600000056", 
4915=>X"00000056000000560000005600000056", 4916=>X"00000056000000560000005600000056", 4917=>X"00000056000000560000005600000056", 4918=>X"00000056000000560000005600000056", 4919=>X"00000056000000560000005600000056", 
4920=>X"00000056000000560000005600000056", 4921=>X"00000056000000560000005600000056", 4922=>X"00000056000000560000005600000056", 4923=>X"00000056000000560000005600000056", 4924=>X"00000056000000560000005600000056", 
4925=>X"00000056000000560000005600000056", 4926=>X"00000056000000560000005600000056", 4927=>X"00000056000000560000005600000056", 4928=>X"00000056000000560000005600000056", 4929=>X"00000056000000560000005600000056", 
4930=>X"00000056000000560000005600000056", 4931=>X"00000056000000560000005600000056", 4932=>X"00000056000000560000005600000056", 4933=>X"00000056000000560000005600000056", 4934=>X"00000056000000560000005600000056", 
4935=>X"00000056000000560000005600000056", 4936=>X"00000055000000550000005500000055", 4937=>X"00000055000000550000005500000055", 4938=>X"00000055000000550000005500000055", 4939=>X"00000055000000550000005500000055", 
4940=>X"00000055000000550000005500000055", 4941=>X"00000055000000550000005500000055", 4942=>X"00000055000000550000005500000055", 4943=>X"00000055000000550000005500000055", 4944=>X"00000055000000550000005500000055", 
4945=>X"00000055000000550000005500000055", 4946=>X"00000055000000550000005500000055", 4947=>X"00000055000000550000005500000055", 4948=>X"00000055000000550000005500000055", 4949=>X"00000055000000550000005500000055", 
4950=>X"00000055000000550000005500000055", 4951=>X"00000055000000550000005500000055", 4952=>X"00000055000000550000005500000055", 4953=>X"00000055000000550000005500000055", 4954=>X"00000055000000550000005500000055", 
4955=>X"00000055000000550000005500000055", 4956=>X"00000055000000550000005500000055", 4957=>X"00000055000000550000005500000055", 4958=>X"00000055000000550000005500000055", 4959=>X"00000055000000550000005500000055", 
4960=>X"00000055000000550000005500000055", 4961=>X"00000055000000550000005500000055", 4962=>X"00000055000000550000005500000055", 4963=>X"00000055000000550000005500000055", 4964=>X"00000055000000550000005500000055", 
4965=>X"00000055000000550000005500000055", 4966=>X"00000055000000550000005500000055", 4967=>X"00000055000000550000005500000055", 4968=>X"00000055000000550000005500000055", 4969=>X"00000055000000550000005500000055", 
4970=>X"00000055000000550000005500000055", 4971=>X"00000055000000550000005500000055", 4972=>X"00000054000000540000005400000055", 4973=>X"00000054000000540000005400000054", 4974=>X"00000054000000540000005400000054", 
4975=>X"00000054000000540000005400000054", 4976=>X"00000054000000540000005400000054", 4977=>X"00000054000000540000005400000054", 4978=>X"00000054000000540000005400000054", 4979=>X"00000054000000540000005400000054", 
4980=>X"00000054000000540000005400000054", 4981=>X"00000054000000540000005400000054", 4982=>X"00000054000000540000005400000054", 4983=>X"00000054000000540000005400000054", 4984=>X"00000054000000540000005400000054", 
4985=>X"00000054000000540000005400000054", 4986=>X"00000054000000540000005400000054", 4987=>X"00000054000000540000005400000054", 4988=>X"00000054000000540000005400000054", 4989=>X"00000054000000540000005400000054", 
4990=>X"00000054000000540000005400000054", 4991=>X"00000054000000540000005400000054", 4992=>X"00000054000000540000005400000054", 4993=>X"00000054000000540000005400000054", 4994=>X"00000054000000540000005400000054", 
4995=>X"00000054000000540000005400000054", 4996=>X"00000054000000540000005400000054", 4997=>X"00000054000000540000005400000054", 4998=>X"00000054000000540000005400000054", 4999=>X"00000054000000540000005400000054", 
5000=>X"00000054000000540000005400000054", 5001=>X"00000054000000540000005400000054", 5002=>X"00000054000000540000005400000054", 5003=>X"00000054000000540000005400000054", 5004=>X"00000054000000540000005400000054", 
5005=>X"00000054000000540000005400000054", 5006=>X"00000054000000540000005400000054", 5007=>X"00000054000000540000005400000054", 5008=>X"00000054000000540000005400000054", 5009=>X"00000053000000530000005300000054", 
5010=>X"00000053000000530000005300000053", 5011=>X"00000053000000530000005300000053", 5012=>X"00000053000000530000005300000053", 5013=>X"00000053000000530000005300000053", 5014=>X"00000053000000530000005300000053", 
5015=>X"00000053000000530000005300000053", 5016=>X"00000053000000530000005300000053", 5017=>X"00000053000000530000005300000053", 5018=>X"00000053000000530000005300000053", 5019=>X"00000053000000530000005300000053", 
5020=>X"00000053000000530000005300000053", 5021=>X"00000053000000530000005300000053", 5022=>X"00000053000000530000005300000053", 5023=>X"00000053000000530000005300000053", 5024=>X"00000053000000530000005300000053", 
5025=>X"00000053000000530000005300000053", 5026=>X"00000053000000530000005300000053", 5027=>X"00000053000000530000005300000053", 5028=>X"00000053000000530000005300000053", 5029=>X"00000053000000530000005300000053", 
5030=>X"00000053000000530000005300000053", 5031=>X"00000053000000530000005300000053", 5032=>X"00000053000000530000005300000053", 5033=>X"00000053000000530000005300000053", 5034=>X"00000053000000530000005300000053", 
5035=>X"00000053000000530000005300000053", 5036=>X"00000053000000530000005300000053", 5037=>X"00000053000000530000005300000053", 5038=>X"00000053000000530000005300000053", 5039=>X"00000053000000530000005300000053", 
5040=>X"00000053000000530000005300000053", 5041=>X"00000053000000530000005300000053", 5042=>X"00000053000000530000005300000053", 5043=>X"00000053000000530000005300000053", 5044=>X"00000053000000530000005300000053", 
5045=>X"00000053000000530000005300000053", 5046=>X"00000053000000530000005300000053", 5047=>X"00000052000000520000005300000053", 5048=>X"00000052000000520000005200000052", 5049=>X"00000052000000520000005200000052", 
5050=>X"00000052000000520000005200000052", 5051=>X"00000052000000520000005200000052", 5052=>X"00000052000000520000005200000052", 5053=>X"00000052000000520000005200000052", 5054=>X"00000052000000520000005200000052", 
5055=>X"00000052000000520000005200000052", 5056=>X"00000052000000520000005200000052", 5057=>X"00000052000000520000005200000052", 5058=>X"00000052000000520000005200000052", 5059=>X"00000052000000520000005200000052", 
5060=>X"00000052000000520000005200000052", 5061=>X"00000052000000520000005200000052", 5062=>X"00000052000000520000005200000052", 5063=>X"00000052000000520000005200000052", 5064=>X"00000052000000520000005200000052", 
5065=>X"00000052000000520000005200000052", 5066=>X"00000052000000520000005200000052", 5067=>X"00000052000000520000005200000052", 5068=>X"00000052000000520000005200000052", 5069=>X"00000052000000520000005200000052", 
5070=>X"00000052000000520000005200000052", 5071=>X"00000052000000520000005200000052", 5072=>X"00000052000000520000005200000052", 5073=>X"00000052000000520000005200000052", 5074=>X"00000052000000520000005200000052", 
5075=>X"00000052000000520000005200000052", 5076=>X"00000052000000520000005200000052", 5077=>X"00000052000000520000005200000052", 5078=>X"00000052000000520000005200000052", 5079=>X"00000052000000520000005200000052", 
5080=>X"00000052000000520000005200000052", 5081=>X"00000052000000520000005200000052", 5082=>X"00000052000000520000005200000052", 5083=>X"00000052000000520000005200000052", 5084=>X"00000052000000520000005200000052", 
5085=>X"00000052000000520000005200000052", 5086=>X"00000051000000510000005100000052", 5087=>X"00000051000000510000005100000051", 5088=>X"00000051000000510000005100000051", 5089=>X"00000051000000510000005100000051", 
5090=>X"00000051000000510000005100000051", 5091=>X"00000051000000510000005100000051", 5092=>X"00000051000000510000005100000051", 5093=>X"00000051000000510000005100000051", 5094=>X"00000051000000510000005100000051", 
5095=>X"00000051000000510000005100000051", 5096=>X"00000051000000510000005100000051", 5097=>X"00000051000000510000005100000051", 5098=>X"00000051000000510000005100000051", 5099=>X"00000051000000510000005100000051", 
5100=>X"00000051000000510000005100000051", 5101=>X"00000051000000510000005100000051", 5102=>X"00000051000000510000005100000051", 5103=>X"00000051000000510000005100000051", 5104=>X"00000051000000510000005100000051", 
5105=>X"00000051000000510000005100000051", 5106=>X"00000051000000510000005100000051", 5107=>X"00000051000000510000005100000051", 5108=>X"00000051000000510000005100000051", 5109=>X"00000051000000510000005100000051", 
5110=>X"00000051000000510000005100000051", 5111=>X"00000051000000510000005100000051", 5112=>X"00000051000000510000005100000051", 5113=>X"00000051000000510000005100000051", 5114=>X"00000051000000510000005100000051", 
5115=>X"00000051000000510000005100000051", 5116=>X"00000051000000510000005100000051", 5117=>X"00000051000000510000005100000051", 5118=>X"00000051000000510000005100000051", 5119=>X"00000051000000510000005100000051", 
5120=>X"00000051000000510000005100000051", 5121=>X"00000051000000510000005100000051", 5122=>X"00000051000000510000005100000051", 5123=>X"00000051000000510000005100000051", 5124=>X"00000051000000510000005100000051", 
5125=>X"00000051000000510000005100000051", 5126=>X"00000050000000500000005000000051", 5127=>X"00000050000000500000005000000050", 5128=>X"00000050000000500000005000000050", 5129=>X"00000050000000500000005000000050", 
5130=>X"00000050000000500000005000000050", 5131=>X"00000050000000500000005000000050", 5132=>X"00000050000000500000005000000050", 5133=>X"00000050000000500000005000000050", 5134=>X"00000050000000500000005000000050", 
5135=>X"00000050000000500000005000000050", 5136=>X"00000050000000500000005000000050", 5137=>X"00000050000000500000005000000050", 5138=>X"00000050000000500000005000000050", 5139=>X"00000050000000500000005000000050", 
5140=>X"00000050000000500000005000000050", 5141=>X"00000050000000500000005000000050", 5142=>X"00000050000000500000005000000050", 5143=>X"00000050000000500000005000000050", 5144=>X"00000050000000500000005000000050", 
5145=>X"00000050000000500000005000000050", 5146=>X"00000050000000500000005000000050", 5147=>X"00000050000000500000005000000050", 5148=>X"00000050000000500000005000000050", 5149=>X"00000050000000500000005000000050", 
5150=>X"00000050000000500000005000000050", 5151=>X"00000050000000500000005000000050", 5152=>X"00000050000000500000005000000050", 5153=>X"00000050000000500000005000000050", 5154=>X"00000050000000500000005000000050", 
5155=>X"00000050000000500000005000000050", 5156=>X"00000050000000500000005000000050", 5157=>X"00000050000000500000005000000050", 5158=>X"00000050000000500000005000000050", 5159=>X"00000050000000500000005000000050", 
5160=>X"00000050000000500000005000000050", 5161=>X"00000050000000500000005000000050", 5162=>X"00000050000000500000005000000050", 5163=>X"00000050000000500000005000000050", 5164=>X"00000050000000500000005000000050", 
5165=>X"00000050000000500000005000000050", 5166=>X"00000050000000500000005000000050", 5167=>X"0000004f0000004f0000004f00000050", 5168=>X"0000004f0000004f0000004f0000004f", 5169=>X"0000004f0000004f0000004f0000004f", 
5170=>X"0000004f0000004f0000004f0000004f", 5171=>X"0000004f0000004f0000004f0000004f", 5172=>X"0000004f0000004f0000004f0000004f", 5173=>X"0000004f0000004f0000004f0000004f", 5174=>X"0000004f0000004f0000004f0000004f", 
5175=>X"0000004f0000004f0000004f0000004f", 5176=>X"0000004f0000004f0000004f0000004f", 5177=>X"0000004f0000004f0000004f0000004f", 5178=>X"0000004f0000004f0000004f0000004f", 5179=>X"0000004f0000004f0000004f0000004f", 
5180=>X"0000004f0000004f0000004f0000004f", 5181=>X"0000004f0000004f0000004f0000004f", 5182=>X"0000004f0000004f0000004f0000004f", 5183=>X"0000004f0000004f0000004f0000004f", 5184=>X"0000004f0000004f0000004f0000004f", 
5185=>X"0000004f0000004f0000004f0000004f", 5186=>X"0000004f0000004f0000004f0000004f", 5187=>X"0000004f0000004f0000004f0000004f", 5188=>X"0000004f0000004f0000004f0000004f", 5189=>X"0000004f0000004f0000004f0000004f", 
5190=>X"0000004f0000004f0000004f0000004f", 5191=>X"0000004f0000004f0000004f0000004f", 5192=>X"0000004f0000004f0000004f0000004f", 5193=>X"0000004f0000004f0000004f0000004f", 5194=>X"0000004f0000004f0000004f0000004f", 
5195=>X"0000004f0000004f0000004f0000004f", 5196=>X"0000004f0000004f0000004f0000004f", 5197=>X"0000004f0000004f0000004f0000004f", 5198=>X"0000004f0000004f0000004f0000004f", 5199=>X"0000004f0000004f0000004f0000004f", 
5200=>X"0000004f0000004f0000004f0000004f", 5201=>X"0000004f0000004f0000004f0000004f", 5202=>X"0000004f0000004f0000004f0000004f", 5203=>X"0000004f0000004f0000004f0000004f", 5204=>X"0000004f0000004f0000004f0000004f", 
5205=>X"0000004f0000004f0000004f0000004f", 5206=>X"0000004f0000004f0000004f0000004f", 5207=>X"0000004f0000004f0000004f0000004f", 5208=>X"0000004f0000004f0000004f0000004f", 5209=>X"0000004e0000004e0000004e0000004f", 
5210=>X"0000004e0000004e0000004e0000004e", 5211=>X"0000004e0000004e0000004e0000004e", 5212=>X"0000004e0000004e0000004e0000004e", 5213=>X"0000004e0000004e0000004e0000004e", 5214=>X"0000004e0000004e0000004e0000004e", 
5215=>X"0000004e0000004e0000004e0000004e", 5216=>X"0000004e0000004e0000004e0000004e", 5217=>X"0000004e0000004e0000004e0000004e", 5218=>X"0000004e0000004e0000004e0000004e", 5219=>X"0000004e0000004e0000004e0000004e", 
5220=>X"0000004e0000004e0000004e0000004e", 5221=>X"0000004e0000004e0000004e0000004e", 5222=>X"0000004e0000004e0000004e0000004e", 5223=>X"0000004e0000004e0000004e0000004e", 5224=>X"0000004e0000004e0000004e0000004e", 
5225=>X"0000004e0000004e0000004e0000004e", 5226=>X"0000004e0000004e0000004e0000004e", 5227=>X"0000004e0000004e0000004e0000004e", 5228=>X"0000004e0000004e0000004e0000004e", 5229=>X"0000004e0000004e0000004e0000004e", 
5230=>X"0000004e0000004e0000004e0000004e", 5231=>X"0000004e0000004e0000004e0000004e", 5232=>X"0000004e0000004e0000004e0000004e", 5233=>X"0000004e0000004e0000004e0000004e", 5234=>X"0000004e0000004e0000004e0000004e", 
5235=>X"0000004e0000004e0000004e0000004e", 5236=>X"0000004e0000004e0000004e0000004e", 5237=>X"0000004e0000004e0000004e0000004e", 5238=>X"0000004e0000004e0000004e0000004e", 5239=>X"0000004e0000004e0000004e0000004e", 
5240=>X"0000004e0000004e0000004e0000004e", 5241=>X"0000004e0000004e0000004e0000004e", 5242=>X"0000004e0000004e0000004e0000004e", 5243=>X"0000004e0000004e0000004e0000004e", 5244=>X"0000004e0000004e0000004e0000004e", 
5245=>X"0000004e0000004e0000004e0000004e", 5246=>X"0000004e0000004e0000004e0000004e", 5247=>X"0000004e0000004e0000004e0000004e", 5248=>X"0000004e0000004e0000004e0000004e", 5249=>X"0000004e0000004e0000004e0000004e", 
5250=>X"0000004e0000004e0000004e0000004e", 5251=>X"0000004e0000004e0000004e0000004e", 5252=>X"0000004d0000004d0000004e0000004e", 5253=>X"0000004d0000004d0000004d0000004d", 5254=>X"0000004d0000004d0000004d0000004d", 
5255=>X"0000004d0000004d0000004d0000004d", 5256=>X"0000004d0000004d0000004d0000004d", 5257=>X"0000004d0000004d0000004d0000004d", 5258=>X"0000004d0000004d0000004d0000004d", 5259=>X"0000004d0000004d0000004d0000004d", 
5260=>X"0000004d0000004d0000004d0000004d", 5261=>X"0000004d0000004d0000004d0000004d", 5262=>X"0000004d0000004d0000004d0000004d", 5263=>X"0000004d0000004d0000004d0000004d", 5264=>X"0000004d0000004d0000004d0000004d", 
5265=>X"0000004d0000004d0000004d0000004d", 5266=>X"0000004d0000004d0000004d0000004d", 5267=>X"0000004d0000004d0000004d0000004d", 5268=>X"0000004d0000004d0000004d0000004d", 5269=>X"0000004d0000004d0000004d0000004d", 
5270=>X"0000004d0000004d0000004d0000004d", 5271=>X"0000004d0000004d0000004d0000004d", 5272=>X"0000004d0000004d0000004d0000004d", 5273=>X"0000004d0000004d0000004d0000004d", 5274=>X"0000004d0000004d0000004d0000004d", 
5275=>X"0000004d0000004d0000004d0000004d", 5276=>X"0000004d0000004d0000004d0000004d", 5277=>X"0000004d0000004d0000004d0000004d", 5278=>X"0000004d0000004d0000004d0000004d", 5279=>X"0000004d0000004d0000004d0000004d", 
5280=>X"0000004d0000004d0000004d0000004d", 5281=>X"0000004d0000004d0000004d0000004d", 5282=>X"0000004d0000004d0000004d0000004d", 5283=>X"0000004d0000004d0000004d0000004d", 5284=>X"0000004d0000004d0000004d0000004d", 
5285=>X"0000004d0000004d0000004d0000004d", 5286=>X"0000004d0000004d0000004d0000004d", 5287=>X"0000004d0000004d0000004d0000004d", 5288=>X"0000004d0000004d0000004d0000004d", 5289=>X"0000004d0000004d0000004d0000004d", 
5290=>X"0000004d0000004d0000004d0000004d", 5291=>X"0000004d0000004d0000004d0000004d", 5292=>X"0000004d0000004d0000004d0000004d", 5293=>X"0000004d0000004d0000004d0000004d", 5294=>X"0000004d0000004d0000004d0000004d", 
5295=>X"0000004d0000004d0000004d0000004d", 5296=>X"0000004c0000004c0000004d0000004d", 5297=>X"0000004c0000004c0000004c0000004c", 5298=>X"0000004c0000004c0000004c0000004c", 5299=>X"0000004c0000004c0000004c0000004c", 
5300=>X"0000004c0000004c0000004c0000004c", 5301=>X"0000004c0000004c0000004c0000004c", 5302=>X"0000004c0000004c0000004c0000004c", 5303=>X"0000004c0000004c0000004c0000004c", 5304=>X"0000004c0000004c0000004c0000004c", 
5305=>X"0000004c0000004c0000004c0000004c", 5306=>X"0000004c0000004c0000004c0000004c", 5307=>X"0000004c0000004c0000004c0000004c", 5308=>X"0000004c0000004c0000004c0000004c", 5309=>X"0000004c0000004c0000004c0000004c", 
5310=>X"0000004c0000004c0000004c0000004c", 5311=>X"0000004c0000004c0000004c0000004c", 5312=>X"0000004c0000004c0000004c0000004c", 5313=>X"0000004c0000004c0000004c0000004c", 5314=>X"0000004c0000004c0000004c0000004c", 
5315=>X"0000004c0000004c0000004c0000004c", 5316=>X"0000004c0000004c0000004c0000004c", 5317=>X"0000004c0000004c0000004c0000004c", 5318=>X"0000004c0000004c0000004c0000004c", 5319=>X"0000004c0000004c0000004c0000004c", 
5320=>X"0000004c0000004c0000004c0000004c", 5321=>X"0000004c0000004c0000004c0000004c", 5322=>X"0000004c0000004c0000004c0000004c", 5323=>X"0000004c0000004c0000004c0000004c", 5324=>X"0000004c0000004c0000004c0000004c", 
5325=>X"0000004c0000004c0000004c0000004c", 5326=>X"0000004c0000004c0000004c0000004c", 5327=>X"0000004c0000004c0000004c0000004c", 5328=>X"0000004c0000004c0000004c0000004c", 5329=>X"0000004c0000004c0000004c0000004c", 
5330=>X"0000004c0000004c0000004c0000004c", 5331=>X"0000004c0000004c0000004c0000004c", 5332=>X"0000004c0000004c0000004c0000004c", 5333=>X"0000004c0000004c0000004c0000004c", 5334=>X"0000004c0000004c0000004c0000004c", 
5335=>X"0000004c0000004c0000004c0000004c", 5336=>X"0000004c0000004c0000004c0000004c", 5337=>X"0000004c0000004c0000004c0000004c", 5338=>X"0000004c0000004c0000004c0000004c", 5339=>X"0000004c0000004c0000004c0000004c", 
5340=>X"0000004c0000004c0000004c0000004c", 5341=>X"0000004c0000004c0000004c0000004c", 5342=>X"0000004b0000004b0000004b0000004b", 5343=>X"0000004b0000004b0000004b0000004b", 5344=>X"0000004b0000004b0000004b0000004b", 
5345=>X"0000004b0000004b0000004b0000004b", 5346=>X"0000004b0000004b0000004b0000004b", 5347=>X"0000004b0000004b0000004b0000004b", 5348=>X"0000004b0000004b0000004b0000004b", 5349=>X"0000004b0000004b0000004b0000004b", 
5350=>X"0000004b0000004b0000004b0000004b", 5351=>X"0000004b0000004b0000004b0000004b", 5352=>X"0000004b0000004b0000004b0000004b", 5353=>X"0000004b0000004b0000004b0000004b", 5354=>X"0000004b0000004b0000004b0000004b", 
5355=>X"0000004b0000004b0000004b0000004b", 5356=>X"0000004b0000004b0000004b0000004b", 5357=>X"0000004b0000004b0000004b0000004b", 5358=>X"0000004b0000004b0000004b0000004b", 5359=>X"0000004b0000004b0000004b0000004b", 
5360=>X"0000004b0000004b0000004b0000004b", 5361=>X"0000004b0000004b0000004b0000004b", 5362=>X"0000004b0000004b0000004b0000004b", 5363=>X"0000004b0000004b0000004b0000004b", 5364=>X"0000004b0000004b0000004b0000004b", 
5365=>X"0000004b0000004b0000004b0000004b", 5366=>X"0000004b0000004b0000004b0000004b", 5367=>X"0000004b0000004b0000004b0000004b", 5368=>X"0000004b0000004b0000004b0000004b", 5369=>X"0000004b0000004b0000004b0000004b", 
5370=>X"0000004b0000004b0000004b0000004b", 5371=>X"0000004b0000004b0000004b0000004b", 5372=>X"0000004b0000004b0000004b0000004b", 5373=>X"0000004b0000004b0000004b0000004b", 5374=>X"0000004b0000004b0000004b0000004b", 
5375=>X"0000004b0000004b0000004b0000004b", 5376=>X"0000004b0000004b0000004b0000004b", 5377=>X"0000004b0000004b0000004b0000004b", 5378=>X"0000004b0000004b0000004b0000004b", 5379=>X"0000004b0000004b0000004b0000004b", 
5380=>X"0000004b0000004b0000004b0000004b", 5381=>X"0000004b0000004b0000004b0000004b", 5382=>X"0000004b0000004b0000004b0000004b", 5383=>X"0000004b0000004b0000004b0000004b", 5384=>X"0000004b0000004b0000004b0000004b", 
5385=>X"0000004b0000004b0000004b0000004b", 5386=>X"0000004b0000004b0000004b0000004b", 5387=>X"0000004b0000004b0000004b0000004b", 5388=>X"0000004a0000004a0000004b0000004b", 5389=>X"0000004a0000004a0000004a0000004a", 
5390=>X"0000004a0000004a0000004a0000004a", 5391=>X"0000004a0000004a0000004a0000004a", 5392=>X"0000004a0000004a0000004a0000004a", 5393=>X"0000004a0000004a0000004a0000004a", 5394=>X"0000004a0000004a0000004a0000004a", 
5395=>X"0000004a0000004a0000004a0000004a", 5396=>X"0000004a0000004a0000004a0000004a", 5397=>X"0000004a0000004a0000004a0000004a", 5398=>X"0000004a0000004a0000004a0000004a", 5399=>X"0000004a0000004a0000004a0000004a", 
5400=>X"0000004a0000004a0000004a0000004a", 5401=>X"0000004a0000004a0000004a0000004a", 5402=>X"0000004a0000004a0000004a0000004a", 5403=>X"0000004a0000004a0000004a0000004a", 5404=>X"0000004a0000004a0000004a0000004a", 
5405=>X"0000004a0000004a0000004a0000004a", 5406=>X"0000004a0000004a0000004a0000004a", 5407=>X"0000004a0000004a0000004a0000004a", 5408=>X"0000004a0000004a0000004a0000004a", 5409=>X"0000004a0000004a0000004a0000004a", 
5410=>X"0000004a0000004a0000004a0000004a", 5411=>X"0000004a0000004a0000004a0000004a", 5412=>X"0000004a0000004a0000004a0000004a", 5413=>X"0000004a0000004a0000004a0000004a", 5414=>X"0000004a0000004a0000004a0000004a", 
5415=>X"0000004a0000004a0000004a0000004a", 5416=>X"0000004a0000004a0000004a0000004a", 5417=>X"0000004a0000004a0000004a0000004a", 5418=>X"0000004a0000004a0000004a0000004a", 5419=>X"0000004a0000004a0000004a0000004a", 
5420=>X"0000004a0000004a0000004a0000004a", 5421=>X"0000004a0000004a0000004a0000004a", 5422=>X"0000004a0000004a0000004a0000004a", 5423=>X"0000004a0000004a0000004a0000004a", 5424=>X"0000004a0000004a0000004a0000004a", 
5425=>X"0000004a0000004a0000004a0000004a", 5426=>X"0000004a0000004a0000004a0000004a", 5427=>X"0000004a0000004a0000004a0000004a", 5428=>X"0000004a0000004a0000004a0000004a", 5429=>X"0000004a0000004a0000004a0000004a", 
5430=>X"0000004a0000004a0000004a0000004a", 5431=>X"0000004a0000004a0000004a0000004a", 5432=>X"0000004a0000004a0000004a0000004a", 5433=>X"0000004a0000004a0000004a0000004a", 5434=>X"0000004a0000004a0000004a0000004a", 
5435=>X"0000004a0000004a0000004a0000004a", 5436=>X"00000049000000490000004a0000004a", 5437=>X"00000049000000490000004900000049", 5438=>X"00000049000000490000004900000049", 5439=>X"00000049000000490000004900000049", 
5440=>X"00000049000000490000004900000049", 5441=>X"00000049000000490000004900000049", 5442=>X"00000049000000490000004900000049", 5443=>X"00000049000000490000004900000049", 5444=>X"00000049000000490000004900000049", 
5445=>X"00000049000000490000004900000049", 5446=>X"00000049000000490000004900000049", 5447=>X"00000049000000490000004900000049", 5448=>X"00000049000000490000004900000049", 5449=>X"00000049000000490000004900000049", 
5450=>X"00000049000000490000004900000049", 5451=>X"00000049000000490000004900000049", 5452=>X"00000049000000490000004900000049", 5453=>X"00000049000000490000004900000049", 5454=>X"00000049000000490000004900000049", 
5455=>X"00000049000000490000004900000049", 5456=>X"00000049000000490000004900000049", 5457=>X"00000049000000490000004900000049", 5458=>X"00000049000000490000004900000049", 5459=>X"00000049000000490000004900000049", 
5460=>X"00000049000000490000004900000049", 5461=>X"00000049000000490000004900000049", 5462=>X"00000049000000490000004900000049", 5463=>X"00000049000000490000004900000049", 5464=>X"00000049000000490000004900000049", 
5465=>X"00000049000000490000004900000049", 5466=>X"00000049000000490000004900000049", 5467=>X"00000049000000490000004900000049", 5468=>X"00000049000000490000004900000049", 5469=>X"00000049000000490000004900000049", 
5470=>X"00000049000000490000004900000049", 5471=>X"00000049000000490000004900000049", 5472=>X"00000049000000490000004900000049", 5473=>X"00000049000000490000004900000049", 5474=>X"00000049000000490000004900000049", 
5475=>X"00000049000000490000004900000049", 5476=>X"00000049000000490000004900000049", 5477=>X"00000049000000490000004900000049", 5478=>X"00000049000000490000004900000049", 5479=>X"00000049000000490000004900000049", 
5480=>X"00000049000000490000004900000049", 5481=>X"00000049000000490000004900000049", 5482=>X"00000049000000490000004900000049", 5483=>X"00000049000000490000004900000049", 5484=>X"00000049000000490000004900000049", 
5485=>X"00000048000000490000004900000049", 5486=>X"00000048000000480000004800000048", 5487=>X"00000048000000480000004800000048", 5488=>X"00000048000000480000004800000048", 5489=>X"00000048000000480000004800000048", 
5490=>X"00000048000000480000004800000048", 5491=>X"00000048000000480000004800000048", 5492=>X"00000048000000480000004800000048", 5493=>X"00000048000000480000004800000048", 5494=>X"00000048000000480000004800000048", 
5495=>X"00000048000000480000004800000048", 5496=>X"00000048000000480000004800000048", 5497=>X"00000048000000480000004800000048", 5498=>X"00000048000000480000004800000048", 5499=>X"00000048000000480000004800000048", 
5500=>X"00000048000000480000004800000048", 5501=>X"00000048000000480000004800000048", 5502=>X"00000048000000480000004800000048", 5503=>X"00000048000000480000004800000048", 5504=>X"00000048000000480000004800000048", 
5505=>X"00000048000000480000004800000048", 5506=>X"00000048000000480000004800000048", 5507=>X"00000048000000480000004800000048", 5508=>X"00000048000000480000004800000048", 5509=>X"00000048000000480000004800000048", 
5510=>X"00000048000000480000004800000048", 5511=>X"00000048000000480000004800000048", 5512=>X"00000048000000480000004800000048", 5513=>X"00000048000000480000004800000048", 5514=>X"00000048000000480000004800000048", 
5515=>X"00000048000000480000004800000048", 5516=>X"00000048000000480000004800000048", 5517=>X"00000048000000480000004800000048", 5518=>X"00000048000000480000004800000048", 5519=>X"00000048000000480000004800000048", 
5520=>X"00000048000000480000004800000048", 5521=>X"00000048000000480000004800000048", 5522=>X"00000048000000480000004800000048", 5523=>X"00000048000000480000004800000048", 5524=>X"00000048000000480000004800000048", 
5525=>X"00000048000000480000004800000048", 5526=>X"00000048000000480000004800000048", 5527=>X"00000048000000480000004800000048", 5528=>X"00000048000000480000004800000048", 5529=>X"00000048000000480000004800000048", 
5530=>X"00000048000000480000004800000048", 5531=>X"00000048000000480000004800000048", 5532=>X"00000048000000480000004800000048", 5533=>X"00000048000000480000004800000048", 5534=>X"00000048000000480000004800000048", 
5535=>X"00000048000000480000004800000048", 5536=>X"00000047000000470000004700000048", 5537=>X"00000047000000470000004700000047", 5538=>X"00000047000000470000004700000047", 5539=>X"00000047000000470000004700000047", 
5540=>X"00000047000000470000004700000047", 5541=>X"00000047000000470000004700000047", 5542=>X"00000047000000470000004700000047", 5543=>X"00000047000000470000004700000047", 5544=>X"00000047000000470000004700000047", 
5545=>X"00000047000000470000004700000047", 5546=>X"00000047000000470000004700000047", 5547=>X"00000047000000470000004700000047", 5548=>X"00000047000000470000004700000047", 5549=>X"00000047000000470000004700000047", 
5550=>X"00000047000000470000004700000047", 5551=>X"00000047000000470000004700000047", 5552=>X"00000047000000470000004700000047", 5553=>X"00000047000000470000004700000047", 5554=>X"00000047000000470000004700000047", 
5555=>X"00000047000000470000004700000047", 5556=>X"00000047000000470000004700000047", 5557=>X"00000047000000470000004700000047", 5558=>X"00000047000000470000004700000047", 5559=>X"00000047000000470000004700000047", 
5560=>X"00000047000000470000004700000047", 5561=>X"00000047000000470000004700000047", 5562=>X"00000047000000470000004700000047", 5563=>X"00000047000000470000004700000047", 5564=>X"00000047000000470000004700000047", 
5565=>X"00000047000000470000004700000047", 5566=>X"00000047000000470000004700000047", 5567=>X"00000047000000470000004700000047", 5568=>X"00000047000000470000004700000047", 5569=>X"00000047000000470000004700000047", 
5570=>X"00000047000000470000004700000047", 5571=>X"00000047000000470000004700000047", 5572=>X"00000047000000470000004700000047", 5573=>X"00000047000000470000004700000047", 5574=>X"00000047000000470000004700000047", 
5575=>X"00000047000000470000004700000047", 5576=>X"00000047000000470000004700000047", 5577=>X"00000047000000470000004700000047", 5578=>X"00000047000000470000004700000047", 5579=>X"00000047000000470000004700000047", 
5580=>X"00000047000000470000004700000047", 5581=>X"00000047000000470000004700000047", 5582=>X"00000047000000470000004700000047", 5583=>X"00000047000000470000004700000047", 5584=>X"00000047000000470000004700000047", 
5585=>X"00000047000000470000004700000047", 5586=>X"00000047000000470000004700000047", 5587=>X"00000047000000470000004700000047", 5588=>X"00000046000000460000004600000047", 5589=>X"00000046000000460000004600000046", 
5590=>X"00000046000000460000004600000046", 5591=>X"00000046000000460000004600000046", 5592=>X"00000046000000460000004600000046", 5593=>X"00000046000000460000004600000046", 5594=>X"00000046000000460000004600000046", 
5595=>X"00000046000000460000004600000046", 5596=>X"00000046000000460000004600000046", 5597=>X"00000046000000460000004600000046", 5598=>X"00000046000000460000004600000046", 5599=>X"00000046000000460000004600000046", 
5600=>X"00000046000000460000004600000046", 5601=>X"00000046000000460000004600000046", 5602=>X"00000046000000460000004600000046", 5603=>X"00000046000000460000004600000046", 5604=>X"00000046000000460000004600000046", 
5605=>X"00000046000000460000004600000046", 5606=>X"00000046000000460000004600000046", 5607=>X"00000046000000460000004600000046", 5608=>X"00000046000000460000004600000046", 5609=>X"00000046000000460000004600000046", 
5610=>X"00000046000000460000004600000046", 5611=>X"00000046000000460000004600000046", 5612=>X"00000046000000460000004600000046", 5613=>X"00000046000000460000004600000046", 5614=>X"00000046000000460000004600000046", 
5615=>X"00000046000000460000004600000046", 5616=>X"00000046000000460000004600000046", 5617=>X"00000046000000460000004600000046", 5618=>X"00000046000000460000004600000046", 5619=>X"00000046000000460000004600000046", 
5620=>X"00000046000000460000004600000046", 5621=>X"00000046000000460000004600000046", 5622=>X"00000046000000460000004600000046", 5623=>X"00000046000000460000004600000046", 5624=>X"00000046000000460000004600000046", 
5625=>X"00000046000000460000004600000046", 5626=>X"00000046000000460000004600000046", 5627=>X"00000046000000460000004600000046", 5628=>X"00000046000000460000004600000046", 5629=>X"00000046000000460000004600000046", 
5630=>X"00000046000000460000004600000046", 5631=>X"00000046000000460000004600000046", 5632=>X"00000046000000460000004600000046", 5633=>X"00000046000000460000004600000046", 5634=>X"00000046000000460000004600000046", 
5635=>X"00000046000000460000004600000046", 5636=>X"00000046000000460000004600000046", 5637=>X"00000046000000460000004600000046", 5638=>X"00000046000000460000004600000046", 5639=>X"00000046000000460000004600000046", 
5640=>X"00000046000000460000004600000046", 5641=>X"00000045000000460000004600000046", 5642=>X"00000045000000450000004500000045", 5643=>X"00000045000000450000004500000045", 5644=>X"00000045000000450000004500000045", 
5645=>X"00000045000000450000004500000045", 5646=>X"00000045000000450000004500000045", 5647=>X"00000045000000450000004500000045", 5648=>X"00000045000000450000004500000045", 5649=>X"00000045000000450000004500000045", 
5650=>X"00000045000000450000004500000045", 5651=>X"00000045000000450000004500000045", 5652=>X"00000045000000450000004500000045", 5653=>X"00000045000000450000004500000045", 5654=>X"00000045000000450000004500000045", 
5655=>X"00000045000000450000004500000045", 5656=>X"00000045000000450000004500000045", 5657=>X"00000045000000450000004500000045", 5658=>X"00000045000000450000004500000045", 5659=>X"00000045000000450000004500000045", 
5660=>X"00000045000000450000004500000045", 5661=>X"00000045000000450000004500000045", 5662=>X"00000045000000450000004500000045", 5663=>X"00000045000000450000004500000045", 5664=>X"00000045000000450000004500000045", 
5665=>X"00000045000000450000004500000045", 5666=>X"00000045000000450000004500000045", 5667=>X"00000045000000450000004500000045", 5668=>X"00000045000000450000004500000045", 5669=>X"00000045000000450000004500000045", 
5670=>X"00000045000000450000004500000045", 5671=>X"00000045000000450000004500000045", 5672=>X"00000045000000450000004500000045", 5673=>X"00000045000000450000004500000045", 5674=>X"00000045000000450000004500000045", 
5675=>X"00000045000000450000004500000045", 5676=>X"00000045000000450000004500000045", 5677=>X"00000045000000450000004500000045", 5678=>X"00000045000000450000004500000045", 5679=>X"00000045000000450000004500000045", 
5680=>X"00000045000000450000004500000045", 5681=>X"00000045000000450000004500000045", 5682=>X"00000045000000450000004500000045", 5683=>X"00000045000000450000004500000045", 5684=>X"00000045000000450000004500000045", 
5685=>X"00000045000000450000004500000045", 5686=>X"00000045000000450000004500000045", 5687=>X"00000045000000450000004500000045", 5688=>X"00000045000000450000004500000045", 5689=>X"00000045000000450000004500000045", 
5690=>X"00000045000000450000004500000045", 5691=>X"00000045000000450000004500000045", 5692=>X"00000045000000450000004500000045", 5693=>X"00000045000000450000004500000045", 5694=>X"00000045000000450000004500000045", 
5695=>X"00000045000000450000004500000045", 5696=>X"00000044000000450000004500000045", 5697=>X"00000044000000440000004400000044", 5698=>X"00000044000000440000004400000044", 5699=>X"00000044000000440000004400000044", 
5700=>X"00000044000000440000004400000044", 5701=>X"00000044000000440000004400000044", 5702=>X"00000044000000440000004400000044", 5703=>X"00000044000000440000004400000044", 5704=>X"00000044000000440000004400000044", 
5705=>X"00000044000000440000004400000044", 5706=>X"00000044000000440000004400000044", 5707=>X"00000044000000440000004400000044", 5708=>X"00000044000000440000004400000044", 5709=>X"00000044000000440000004400000044", 
5710=>X"00000044000000440000004400000044", 5711=>X"00000044000000440000004400000044", 5712=>X"00000044000000440000004400000044", 5713=>X"00000044000000440000004400000044", 5714=>X"00000044000000440000004400000044", 
5715=>X"00000044000000440000004400000044", 5716=>X"00000044000000440000004400000044", 5717=>X"00000044000000440000004400000044", 5718=>X"00000044000000440000004400000044", 5719=>X"00000044000000440000004400000044", 
5720=>X"00000044000000440000004400000044", 5721=>X"00000044000000440000004400000044", 5722=>X"00000044000000440000004400000044", 5723=>X"00000044000000440000004400000044", 5724=>X"00000044000000440000004400000044", 
5725=>X"00000044000000440000004400000044", 5726=>X"00000044000000440000004400000044", 5727=>X"00000044000000440000004400000044", 5728=>X"00000044000000440000004400000044", 5729=>X"00000044000000440000004400000044", 
5730=>X"00000044000000440000004400000044", 5731=>X"00000044000000440000004400000044", 5732=>X"00000044000000440000004400000044", 5733=>X"00000044000000440000004400000044", 5734=>X"00000044000000440000004400000044", 
5735=>X"00000044000000440000004400000044", 5736=>X"00000044000000440000004400000044", 5737=>X"00000044000000440000004400000044", 5738=>X"00000044000000440000004400000044", 5739=>X"00000044000000440000004400000044", 
5740=>X"00000044000000440000004400000044", 5741=>X"00000044000000440000004400000044", 5742=>X"00000044000000440000004400000044", 5743=>X"00000044000000440000004400000044", 5744=>X"00000044000000440000004400000044", 
5745=>X"00000044000000440000004400000044", 5746=>X"00000044000000440000004400000044", 5747=>X"00000044000000440000004400000044", 5748=>X"00000044000000440000004400000044", 5749=>X"00000044000000440000004400000044", 
5750=>X"00000044000000440000004400000044", 5751=>X"00000044000000440000004400000044", 5752=>X"00000044000000440000004400000044", 5753=>X"00000043000000430000004400000044", 5754=>X"00000043000000430000004300000043", 
5755=>X"00000043000000430000004300000043", 5756=>X"00000043000000430000004300000043", 5757=>X"00000043000000430000004300000043", 5758=>X"00000043000000430000004300000043", 5759=>X"00000043000000430000004300000043", 
5760=>X"00000043000000430000004300000043", 5761=>X"00000043000000430000004300000043", 5762=>X"00000043000000430000004300000043", 5763=>X"00000043000000430000004300000043", 5764=>X"00000043000000430000004300000043", 
5765=>X"00000043000000430000004300000043", 5766=>X"00000043000000430000004300000043", 5767=>X"00000043000000430000004300000043", 5768=>X"00000043000000430000004300000043", 5769=>X"00000043000000430000004300000043", 
5770=>X"00000043000000430000004300000043", 5771=>X"00000043000000430000004300000043", 5772=>X"00000043000000430000004300000043", 5773=>X"00000043000000430000004300000043", 5774=>X"00000043000000430000004300000043", 
5775=>X"00000043000000430000004300000043", 5776=>X"00000043000000430000004300000043", 5777=>X"00000043000000430000004300000043", 5778=>X"00000043000000430000004300000043", 5779=>X"00000043000000430000004300000043", 
5780=>X"00000043000000430000004300000043", 5781=>X"00000043000000430000004300000043", 5782=>X"00000043000000430000004300000043", 5783=>X"00000043000000430000004300000043", 5784=>X"00000043000000430000004300000043", 
5785=>X"00000043000000430000004300000043", 5786=>X"00000043000000430000004300000043", 5787=>X"00000043000000430000004300000043", 5788=>X"00000043000000430000004300000043", 5789=>X"00000043000000430000004300000043", 
5790=>X"00000043000000430000004300000043", 5791=>X"00000043000000430000004300000043", 5792=>X"00000043000000430000004300000043", 5793=>X"00000043000000430000004300000043", 5794=>X"00000043000000430000004300000043", 
5795=>X"00000043000000430000004300000043", 5796=>X"00000043000000430000004300000043", 5797=>X"00000043000000430000004300000043", 5798=>X"00000043000000430000004300000043", 5799=>X"00000043000000430000004300000043", 
5800=>X"00000043000000430000004300000043", 5801=>X"00000043000000430000004300000043", 5802=>X"00000043000000430000004300000043", 5803=>X"00000043000000430000004300000043", 5804=>X"00000043000000430000004300000043", 
5805=>X"00000043000000430000004300000043", 5806=>X"00000043000000430000004300000043", 5807=>X"00000043000000430000004300000043", 5808=>X"00000043000000430000004300000043", 5809=>X"00000043000000430000004300000043", 
5810=>X"00000043000000430000004300000043", 5811=>X"00000043000000430000004300000043", 5812=>X"00000042000000420000004200000042", 5813=>X"00000042000000420000004200000042", 5814=>X"00000042000000420000004200000042", 
5815=>X"00000042000000420000004200000042", 5816=>X"00000042000000420000004200000042", 5817=>X"00000042000000420000004200000042", 5818=>X"00000042000000420000004200000042", 5819=>X"00000042000000420000004200000042", 
5820=>X"00000042000000420000004200000042", 5821=>X"00000042000000420000004200000042", 5822=>X"00000042000000420000004200000042", 5823=>X"00000042000000420000004200000042", 5824=>X"00000042000000420000004200000042", 
5825=>X"00000042000000420000004200000042", 5826=>X"00000042000000420000004200000042", 5827=>X"00000042000000420000004200000042", 5828=>X"00000042000000420000004200000042", 5829=>X"00000042000000420000004200000042", 
5830=>X"00000042000000420000004200000042", 5831=>X"00000042000000420000004200000042", 5832=>X"00000042000000420000004200000042", 5833=>X"00000042000000420000004200000042", 5834=>X"00000042000000420000004200000042", 
5835=>X"00000042000000420000004200000042", 5836=>X"00000042000000420000004200000042", 5837=>X"00000042000000420000004200000042", 5838=>X"00000042000000420000004200000042", 5839=>X"00000042000000420000004200000042", 
5840=>X"00000042000000420000004200000042", 5841=>X"00000042000000420000004200000042", 5842=>X"00000042000000420000004200000042", 5843=>X"00000042000000420000004200000042", 5844=>X"00000042000000420000004200000042", 
5845=>X"00000042000000420000004200000042", 5846=>X"00000042000000420000004200000042", 5847=>X"00000042000000420000004200000042", 5848=>X"00000042000000420000004200000042", 5849=>X"00000042000000420000004200000042", 
5850=>X"00000042000000420000004200000042", 5851=>X"00000042000000420000004200000042", 5852=>X"00000042000000420000004200000042", 5853=>X"00000042000000420000004200000042", 5854=>X"00000042000000420000004200000042", 
5855=>X"00000042000000420000004200000042", 5856=>X"00000042000000420000004200000042", 5857=>X"00000042000000420000004200000042", 5858=>X"00000042000000420000004200000042", 5859=>X"00000042000000420000004200000042", 
5860=>X"00000042000000420000004200000042", 5861=>X"00000042000000420000004200000042", 5862=>X"00000042000000420000004200000042", 5863=>X"00000042000000420000004200000042", 5864=>X"00000042000000420000004200000042", 
5865=>X"00000042000000420000004200000042", 5866=>X"00000042000000420000004200000042", 5867=>X"00000042000000420000004200000042", 5868=>X"00000042000000420000004200000042", 5869=>X"00000042000000420000004200000042", 
5870=>X"00000042000000420000004200000042", 5871=>X"00000042000000420000004200000042", 5872=>X"00000041000000410000004100000041", 5873=>X"00000041000000410000004100000041", 5874=>X"00000041000000410000004100000041", 
5875=>X"00000041000000410000004100000041", 5876=>X"00000041000000410000004100000041", 5877=>X"00000041000000410000004100000041", 5878=>X"00000041000000410000004100000041", 5879=>X"00000041000000410000004100000041", 
5880=>X"00000041000000410000004100000041", 5881=>X"00000041000000410000004100000041", 5882=>X"00000041000000410000004100000041", 5883=>X"00000041000000410000004100000041", 5884=>X"00000041000000410000004100000041", 
5885=>X"00000041000000410000004100000041", 5886=>X"00000041000000410000004100000041", 5887=>X"00000041000000410000004100000041", 5888=>X"00000041000000410000004100000041", 5889=>X"00000041000000410000004100000041", 
5890=>X"00000041000000410000004100000041", 5891=>X"00000041000000410000004100000041", 5892=>X"00000041000000410000004100000041", 5893=>X"00000041000000410000004100000041", 5894=>X"00000041000000410000004100000041", 
5895=>X"00000041000000410000004100000041", 5896=>X"00000041000000410000004100000041", 5897=>X"00000041000000410000004100000041", 5898=>X"00000041000000410000004100000041", 5899=>X"00000041000000410000004100000041", 
5900=>X"00000041000000410000004100000041", 5901=>X"00000041000000410000004100000041", 5902=>X"00000041000000410000004100000041", 5903=>X"00000041000000410000004100000041", 5904=>X"00000041000000410000004100000041", 
5905=>X"00000041000000410000004100000041", 5906=>X"00000041000000410000004100000041", 5907=>X"00000041000000410000004100000041", 5908=>X"00000041000000410000004100000041", 5909=>X"00000041000000410000004100000041", 
5910=>X"00000041000000410000004100000041", 5911=>X"00000041000000410000004100000041", 5912=>X"00000041000000410000004100000041", 5913=>X"00000041000000410000004100000041", 5914=>X"00000041000000410000004100000041", 
5915=>X"00000041000000410000004100000041", 5916=>X"00000041000000410000004100000041", 5917=>X"00000041000000410000004100000041", 5918=>X"00000041000000410000004100000041", 5919=>X"00000041000000410000004100000041", 
5920=>X"00000041000000410000004100000041", 5921=>X"00000041000000410000004100000041", 5922=>X"00000041000000410000004100000041", 5923=>X"00000041000000410000004100000041", 5924=>X"00000041000000410000004100000041", 
5925=>X"00000041000000410000004100000041", 5926=>X"00000041000000410000004100000041", 5927=>X"00000041000000410000004100000041", 5928=>X"00000041000000410000004100000041", 5929=>X"00000041000000410000004100000041", 
5930=>X"00000041000000410000004100000041", 5931=>X"00000041000000410000004100000041", 5932=>X"00000041000000410000004100000041", 5933=>X"00000041000000410000004100000041", 5934=>X"00000040000000400000004000000040", 
5935=>X"00000040000000400000004000000040", 5936=>X"00000040000000400000004000000040", 5937=>X"00000040000000400000004000000040", 5938=>X"00000040000000400000004000000040", 5939=>X"00000040000000400000004000000040", 
5940=>X"00000040000000400000004000000040", 5941=>X"00000040000000400000004000000040", 5942=>X"00000040000000400000004000000040", 5943=>X"00000040000000400000004000000040", 5944=>X"00000040000000400000004000000040", 
5945=>X"00000040000000400000004000000040", 5946=>X"00000040000000400000004000000040", 5947=>X"00000040000000400000004000000040", 5948=>X"00000040000000400000004000000040", 5949=>X"00000040000000400000004000000040", 
5950=>X"00000040000000400000004000000040", 5951=>X"00000040000000400000004000000040", 5952=>X"00000040000000400000004000000040", 5953=>X"00000040000000400000004000000040", 5954=>X"00000040000000400000004000000040", 
5955=>X"00000040000000400000004000000040", 5956=>X"00000040000000400000004000000040", 5957=>X"00000040000000400000004000000040", 5958=>X"00000040000000400000004000000040", 5959=>X"00000040000000400000004000000040", 
5960=>X"00000040000000400000004000000040", 5961=>X"00000040000000400000004000000040", 5962=>X"00000040000000400000004000000040", 5963=>X"00000040000000400000004000000040", 5964=>X"00000040000000400000004000000040", 
5965=>X"00000040000000400000004000000040", 5966=>X"00000040000000400000004000000040", 5967=>X"00000040000000400000004000000040", 5968=>X"00000040000000400000004000000040", 5969=>X"00000040000000400000004000000040", 
5970=>X"00000040000000400000004000000040", 5971=>X"00000040000000400000004000000040", 5972=>X"00000040000000400000004000000040", 5973=>X"00000040000000400000004000000040", 5974=>X"00000040000000400000004000000040", 
5975=>X"00000040000000400000004000000040", 5976=>X"00000040000000400000004000000040", 5977=>X"00000040000000400000004000000040", 5978=>X"00000040000000400000004000000040", 5979=>X"00000040000000400000004000000040", 
5980=>X"00000040000000400000004000000040", 5981=>X"00000040000000400000004000000040", 5982=>X"00000040000000400000004000000040", 5983=>X"00000040000000400000004000000040", 5984=>X"00000040000000400000004000000040", 
5985=>X"00000040000000400000004000000040", 5986=>X"00000040000000400000004000000040", 5987=>X"00000040000000400000004000000040", 5988=>X"00000040000000400000004000000040", 5989=>X"00000040000000400000004000000040", 
5990=>X"00000040000000400000004000000040", 5991=>X"00000040000000400000004000000040", 5992=>X"00000040000000400000004000000040", 5993=>X"00000040000000400000004000000040", 5994=>X"00000040000000400000004000000040", 
5995=>X"00000040000000400000004000000040", 5996=>X"00000040000000400000004000000040", 5997=>X"00000040000000400000004000000040", 5998=>X"0000003f0000003f0000003f00000040", 5999=>X"0000003f0000003f0000003f0000003f", 
6000=>X"0000003f0000003f0000003f0000003f", 6001=>X"0000003f0000003f0000003f0000003f", 6002=>X"0000003f0000003f0000003f0000003f", 6003=>X"0000003f0000003f0000003f0000003f", 6004=>X"0000003f0000003f0000003f0000003f", 
6005=>X"0000003f0000003f0000003f0000003f", 6006=>X"0000003f0000003f0000003f0000003f", 6007=>X"0000003f0000003f0000003f0000003f", 6008=>X"0000003f0000003f0000003f0000003f", 6009=>X"0000003f0000003f0000003f0000003f", 
6010=>X"0000003f0000003f0000003f0000003f", 6011=>X"0000003f0000003f0000003f0000003f", 6012=>X"0000003f0000003f0000003f0000003f", 6013=>X"0000003f0000003f0000003f0000003f", 6014=>X"0000003f0000003f0000003f0000003f", 
6015=>X"0000003f0000003f0000003f0000003f", 6016=>X"0000003f0000003f0000003f0000003f", 6017=>X"0000003f0000003f0000003f0000003f", 6018=>X"0000003f0000003f0000003f0000003f", 6019=>X"0000003f0000003f0000003f0000003f", 
6020=>X"0000003f0000003f0000003f0000003f", 6021=>X"0000003f0000003f0000003f0000003f", 6022=>X"0000003f0000003f0000003f0000003f", 6023=>X"0000003f0000003f0000003f0000003f", 6024=>X"0000003f0000003f0000003f0000003f", 
6025=>X"0000003f0000003f0000003f0000003f", 6026=>X"0000003f0000003f0000003f0000003f", 6027=>X"0000003f0000003f0000003f0000003f", 6028=>X"0000003f0000003f0000003f0000003f", 6029=>X"0000003f0000003f0000003f0000003f", 
6030=>X"0000003f0000003f0000003f0000003f", 6031=>X"0000003f0000003f0000003f0000003f", 6032=>X"0000003f0000003f0000003f0000003f", 6033=>X"0000003f0000003f0000003f0000003f", 6034=>X"0000003f0000003f0000003f0000003f", 
6035=>X"0000003f0000003f0000003f0000003f", 6036=>X"0000003f0000003f0000003f0000003f", 6037=>X"0000003f0000003f0000003f0000003f", 6038=>X"0000003f0000003f0000003f0000003f", 6039=>X"0000003f0000003f0000003f0000003f", 
6040=>X"0000003f0000003f0000003f0000003f", 6041=>X"0000003f0000003f0000003f0000003f", 6042=>X"0000003f0000003f0000003f0000003f", 6043=>X"0000003f0000003f0000003f0000003f", 6044=>X"0000003f0000003f0000003f0000003f", 
6045=>X"0000003f0000003f0000003f0000003f", 6046=>X"0000003f0000003f0000003f0000003f", 6047=>X"0000003f0000003f0000003f0000003f", 6048=>X"0000003f0000003f0000003f0000003f", 6049=>X"0000003f0000003f0000003f0000003f", 
6050=>X"0000003f0000003f0000003f0000003f", 6051=>X"0000003f0000003f0000003f0000003f", 6052=>X"0000003f0000003f0000003f0000003f", 6053=>X"0000003f0000003f0000003f0000003f", 6054=>X"0000003f0000003f0000003f0000003f", 
6055=>X"0000003f0000003f0000003f0000003f", 6056=>X"0000003f0000003f0000003f0000003f", 6057=>X"0000003f0000003f0000003f0000003f", 6058=>X"0000003f0000003f0000003f0000003f", 6059=>X"0000003f0000003f0000003f0000003f", 
6060=>X"0000003f0000003f0000003f0000003f", 6061=>X"0000003f0000003f0000003f0000003f", 6062=>X"0000003f0000003f0000003f0000003f", 6063=>X"0000003f0000003f0000003f0000003f", 6064=>X"0000003e0000003e0000003e0000003f", 
6065=>X"0000003e0000003e0000003e0000003e", 6066=>X"0000003e0000003e0000003e0000003e", 6067=>X"0000003e0000003e0000003e0000003e", 6068=>X"0000003e0000003e0000003e0000003e", 6069=>X"0000003e0000003e0000003e0000003e", 
6070=>X"0000003e0000003e0000003e0000003e", 6071=>X"0000003e0000003e0000003e0000003e", 6072=>X"0000003e0000003e0000003e0000003e", 6073=>X"0000003e0000003e0000003e0000003e", 6074=>X"0000003e0000003e0000003e0000003e", 
6075=>X"0000003e0000003e0000003e0000003e", 6076=>X"0000003e0000003e0000003e0000003e", 6077=>X"0000003e0000003e0000003e0000003e", 6078=>X"0000003e0000003e0000003e0000003e", 6079=>X"0000003e0000003e0000003e0000003e", 
6080=>X"0000003e0000003e0000003e0000003e", 6081=>X"0000003e0000003e0000003e0000003e", 6082=>X"0000003e0000003e0000003e0000003e", 6083=>X"0000003e0000003e0000003e0000003e", 6084=>X"0000003e0000003e0000003e0000003e", 
6085=>X"0000003e0000003e0000003e0000003e", 6086=>X"0000003e0000003e0000003e0000003e", 6087=>X"0000003e0000003e0000003e0000003e", 6088=>X"0000003e0000003e0000003e0000003e", 6089=>X"0000003e0000003e0000003e0000003e", 
6090=>X"0000003e0000003e0000003e0000003e", 6091=>X"0000003e0000003e0000003e0000003e", 6092=>X"0000003e0000003e0000003e0000003e", 6093=>X"0000003e0000003e0000003e0000003e", 6094=>X"0000003e0000003e0000003e0000003e", 
6095=>X"0000003e0000003e0000003e0000003e", 6096=>X"0000003e0000003e0000003e0000003e", 6097=>X"0000003e0000003e0000003e0000003e", 6098=>X"0000003e0000003e0000003e0000003e", 6099=>X"0000003e0000003e0000003e0000003e", 
6100=>X"0000003e0000003e0000003e0000003e", 6101=>X"0000003e0000003e0000003e0000003e", 6102=>X"0000003e0000003e0000003e0000003e", 6103=>X"0000003e0000003e0000003e0000003e", 6104=>X"0000003e0000003e0000003e0000003e", 
6105=>X"0000003e0000003e0000003e0000003e", 6106=>X"0000003e0000003e0000003e0000003e", 6107=>X"0000003e0000003e0000003e0000003e", 6108=>X"0000003e0000003e0000003e0000003e", 6109=>X"0000003e0000003e0000003e0000003e", 
6110=>X"0000003e0000003e0000003e0000003e", 6111=>X"0000003e0000003e0000003e0000003e", 6112=>X"0000003e0000003e0000003e0000003e", 6113=>X"0000003e0000003e0000003e0000003e", 6114=>X"0000003e0000003e0000003e0000003e", 
6115=>X"0000003e0000003e0000003e0000003e", 6116=>X"0000003e0000003e0000003e0000003e", 6117=>X"0000003e0000003e0000003e0000003e", 6118=>X"0000003e0000003e0000003e0000003e", 6119=>X"0000003e0000003e0000003e0000003e", 
6120=>X"0000003e0000003e0000003e0000003e", 6121=>X"0000003e0000003e0000003e0000003e", 6122=>X"0000003e0000003e0000003e0000003e", 6123=>X"0000003e0000003e0000003e0000003e", 6124=>X"0000003e0000003e0000003e0000003e", 
6125=>X"0000003e0000003e0000003e0000003e", 6126=>X"0000003e0000003e0000003e0000003e", 6127=>X"0000003e0000003e0000003e0000003e", 6128=>X"0000003e0000003e0000003e0000003e", 6129=>X"0000003e0000003e0000003e0000003e", 
6130=>X"0000003e0000003e0000003e0000003e", 6131=>X"0000003e0000003e0000003e0000003e", 6132=>X"0000003d0000003d0000003e0000003e", 6133=>X"0000003d0000003d0000003d0000003d", 6134=>X"0000003d0000003d0000003d0000003d", 
6135=>X"0000003d0000003d0000003d0000003d", 6136=>X"0000003d0000003d0000003d0000003d", 6137=>X"0000003d0000003d0000003d0000003d", 6138=>X"0000003d0000003d0000003d0000003d", 6139=>X"0000003d0000003d0000003d0000003d", 
6140=>X"0000003d0000003d0000003d0000003d", 6141=>X"0000003d0000003d0000003d0000003d", 6142=>X"0000003d0000003d0000003d0000003d", 6143=>X"0000003d0000003d0000003d0000003d", 6144=>X"0000003d0000003d0000003d0000003d", 
6145=>X"0000003d0000003d0000003d0000003d", 6146=>X"0000003d0000003d0000003d0000003d", 6147=>X"0000003d0000003d0000003d0000003d", 6148=>X"0000003d0000003d0000003d0000003d", 6149=>X"0000003d0000003d0000003d0000003d", 
6150=>X"0000003d0000003d0000003d0000003d", 6151=>X"0000003d0000003d0000003d0000003d", 6152=>X"0000003d0000003d0000003d0000003d", 6153=>X"0000003d0000003d0000003d0000003d", 6154=>X"0000003d0000003d0000003d0000003d", 
6155=>X"0000003d0000003d0000003d0000003d", 6156=>X"0000003d0000003d0000003d0000003d", 6157=>X"0000003d0000003d0000003d0000003d", 6158=>X"0000003d0000003d0000003d0000003d", 6159=>X"0000003d0000003d0000003d0000003d", 
6160=>X"0000003d0000003d0000003d0000003d", 6161=>X"0000003d0000003d0000003d0000003d", 6162=>X"0000003d0000003d0000003d0000003d", 6163=>X"0000003d0000003d0000003d0000003d", 6164=>X"0000003d0000003d0000003d0000003d", 
6165=>X"0000003d0000003d0000003d0000003d", 6166=>X"0000003d0000003d0000003d0000003d", 6167=>X"0000003d0000003d0000003d0000003d", 6168=>X"0000003d0000003d0000003d0000003d", 6169=>X"0000003d0000003d0000003d0000003d", 
6170=>X"0000003d0000003d0000003d0000003d", 6171=>X"0000003d0000003d0000003d0000003d", 6172=>X"0000003d0000003d0000003d0000003d", 6173=>X"0000003d0000003d0000003d0000003d", 6174=>X"0000003d0000003d0000003d0000003d", 
6175=>X"0000003d0000003d0000003d0000003d", 6176=>X"0000003d0000003d0000003d0000003d", 6177=>X"0000003d0000003d0000003d0000003d", 6178=>X"0000003d0000003d0000003d0000003d", 6179=>X"0000003d0000003d0000003d0000003d", 
6180=>X"0000003d0000003d0000003d0000003d", 6181=>X"0000003d0000003d0000003d0000003d", 6182=>X"0000003d0000003d0000003d0000003d", 6183=>X"0000003d0000003d0000003d0000003d", 6184=>X"0000003d0000003d0000003d0000003d", 
6185=>X"0000003d0000003d0000003d0000003d", 6186=>X"0000003d0000003d0000003d0000003d", 6187=>X"0000003d0000003d0000003d0000003d", 6188=>X"0000003d0000003d0000003d0000003d", 6189=>X"0000003d0000003d0000003d0000003d", 
6190=>X"0000003d0000003d0000003d0000003d", 6191=>X"0000003d0000003d0000003d0000003d", 6192=>X"0000003d0000003d0000003d0000003d", 6193=>X"0000003d0000003d0000003d0000003d", 6194=>X"0000003d0000003d0000003d0000003d", 
6195=>X"0000003d0000003d0000003d0000003d", 6196=>X"0000003d0000003d0000003d0000003d", 6197=>X"0000003d0000003d0000003d0000003d", 6198=>X"0000003d0000003d0000003d0000003d", 6199=>X"0000003d0000003d0000003d0000003d", 
6200=>X"0000003d0000003d0000003d0000003d", 6201=>X"0000003d0000003d0000003d0000003d", 6202=>X"0000003c0000003d0000003d0000003d", 6203=>X"0000003c0000003c0000003c0000003c", 6204=>X"0000003c0000003c0000003c0000003c", 
6205=>X"0000003c0000003c0000003c0000003c", 6206=>X"0000003c0000003c0000003c0000003c", 6207=>X"0000003c0000003c0000003c0000003c", 6208=>X"0000003c0000003c0000003c0000003c", 6209=>X"0000003c0000003c0000003c0000003c", 
6210=>X"0000003c0000003c0000003c0000003c", 6211=>X"0000003c0000003c0000003c0000003c", 6212=>X"0000003c0000003c0000003c0000003c", 6213=>X"0000003c0000003c0000003c0000003c", 6214=>X"0000003c0000003c0000003c0000003c", 
6215=>X"0000003c0000003c0000003c0000003c", 6216=>X"0000003c0000003c0000003c0000003c", 6217=>X"0000003c0000003c0000003c0000003c", 6218=>X"0000003c0000003c0000003c0000003c", 6219=>X"0000003c0000003c0000003c0000003c", 
6220=>X"0000003c0000003c0000003c0000003c", 6221=>X"0000003c0000003c0000003c0000003c", 6222=>X"0000003c0000003c0000003c0000003c", 6223=>X"0000003c0000003c0000003c0000003c", 6224=>X"0000003c0000003c0000003c0000003c", 
6225=>X"0000003c0000003c0000003c0000003c", 6226=>X"0000003c0000003c0000003c0000003c", 6227=>X"0000003c0000003c0000003c0000003c", 6228=>X"0000003c0000003c0000003c0000003c", 6229=>X"0000003c0000003c0000003c0000003c", 
6230=>X"0000003c0000003c0000003c0000003c", 6231=>X"0000003c0000003c0000003c0000003c", 6232=>X"0000003c0000003c0000003c0000003c", 6233=>X"0000003c0000003c0000003c0000003c", 6234=>X"0000003c0000003c0000003c0000003c", 
6235=>X"0000003c0000003c0000003c0000003c", 6236=>X"0000003c0000003c0000003c0000003c", 6237=>X"0000003c0000003c0000003c0000003c", 6238=>X"0000003c0000003c0000003c0000003c", 6239=>X"0000003c0000003c0000003c0000003c", 
6240=>X"0000003c0000003c0000003c0000003c", 6241=>X"0000003c0000003c0000003c0000003c", 6242=>X"0000003c0000003c0000003c0000003c", 6243=>X"0000003c0000003c0000003c0000003c", 6244=>X"0000003c0000003c0000003c0000003c", 
6245=>X"0000003c0000003c0000003c0000003c", 6246=>X"0000003c0000003c0000003c0000003c", 6247=>X"0000003c0000003c0000003c0000003c", 6248=>X"0000003c0000003c0000003c0000003c", 6249=>X"0000003c0000003c0000003c0000003c", 
6250=>X"0000003c0000003c0000003c0000003c", 6251=>X"0000003c0000003c0000003c0000003c", 6252=>X"0000003c0000003c0000003c0000003c", 6253=>X"0000003c0000003c0000003c0000003c", 6254=>X"0000003c0000003c0000003c0000003c", 
6255=>X"0000003c0000003c0000003c0000003c", 6256=>X"0000003c0000003c0000003c0000003c", 6257=>X"0000003c0000003c0000003c0000003c", 6258=>X"0000003c0000003c0000003c0000003c", 6259=>X"0000003c0000003c0000003c0000003c", 
6260=>X"0000003c0000003c0000003c0000003c", 6261=>X"0000003c0000003c0000003c0000003c", 6262=>X"0000003c0000003c0000003c0000003c", 6263=>X"0000003c0000003c0000003c0000003c", 6264=>X"0000003c0000003c0000003c0000003c", 
6265=>X"0000003c0000003c0000003c0000003c", 6266=>X"0000003c0000003c0000003c0000003c", 6267=>X"0000003c0000003c0000003c0000003c", 6268=>X"0000003c0000003c0000003c0000003c", 6269=>X"0000003c0000003c0000003c0000003c", 
6270=>X"0000003c0000003c0000003c0000003c", 6271=>X"0000003c0000003c0000003c0000003c", 6272=>X"0000003c0000003c0000003c0000003c", 6273=>X"0000003c0000003c0000003c0000003c", 6274=>X"0000003c0000003c0000003c0000003c", 
6275=>X"0000003b0000003c0000003c0000003c", 6276=>X"0000003b0000003b0000003b0000003b", 6277=>X"0000003b0000003b0000003b0000003b", 6278=>X"0000003b0000003b0000003b0000003b", 6279=>X"0000003b0000003b0000003b0000003b", 
6280=>X"0000003b0000003b0000003b0000003b", 6281=>X"0000003b0000003b0000003b0000003b", 6282=>X"0000003b0000003b0000003b0000003b", 6283=>X"0000003b0000003b0000003b0000003b", 6284=>X"0000003b0000003b0000003b0000003b", 
6285=>X"0000003b0000003b0000003b0000003b", 6286=>X"0000003b0000003b0000003b0000003b", 6287=>X"0000003b0000003b0000003b0000003b", 6288=>X"0000003b0000003b0000003b0000003b", 6289=>X"0000003b0000003b0000003b0000003b", 
6290=>X"0000003b0000003b0000003b0000003b", 6291=>X"0000003b0000003b0000003b0000003b", 6292=>X"0000003b0000003b0000003b0000003b", 6293=>X"0000003b0000003b0000003b0000003b", 6294=>X"0000003b0000003b0000003b0000003b", 
6295=>X"0000003b0000003b0000003b0000003b", 6296=>X"0000003b0000003b0000003b0000003b", 6297=>X"0000003b0000003b0000003b0000003b", 6298=>X"0000003b0000003b0000003b0000003b", 6299=>X"0000003b0000003b0000003b0000003b", 
6300=>X"0000003b0000003b0000003b0000003b", 6301=>X"0000003b0000003b0000003b0000003b", 6302=>X"0000003b0000003b0000003b0000003b", 6303=>X"0000003b0000003b0000003b0000003b", 6304=>X"0000003b0000003b0000003b0000003b", 
6305=>X"0000003b0000003b0000003b0000003b", 6306=>X"0000003b0000003b0000003b0000003b", 6307=>X"0000003b0000003b0000003b0000003b", 6308=>X"0000003b0000003b0000003b0000003b", 6309=>X"0000003b0000003b0000003b0000003b", 
6310=>X"0000003b0000003b0000003b0000003b", 6311=>X"0000003b0000003b0000003b0000003b", 6312=>X"0000003b0000003b0000003b0000003b", 6313=>X"0000003b0000003b0000003b0000003b", 6314=>X"0000003b0000003b0000003b0000003b", 
6315=>X"0000003b0000003b0000003b0000003b", 6316=>X"0000003b0000003b0000003b0000003b", 6317=>X"0000003b0000003b0000003b0000003b", 6318=>X"0000003b0000003b0000003b0000003b", 6319=>X"0000003b0000003b0000003b0000003b", 
6320=>X"0000003b0000003b0000003b0000003b", 6321=>X"0000003b0000003b0000003b0000003b", 6322=>X"0000003b0000003b0000003b0000003b", 6323=>X"0000003b0000003b0000003b0000003b", 6324=>X"0000003b0000003b0000003b0000003b", 
6325=>X"0000003b0000003b0000003b0000003b", 6326=>X"0000003b0000003b0000003b0000003b", 6327=>X"0000003b0000003b0000003b0000003b", 6328=>X"0000003b0000003b0000003b0000003b", 6329=>X"0000003b0000003b0000003b0000003b", 
6330=>X"0000003b0000003b0000003b0000003b", 6331=>X"0000003b0000003b0000003b0000003b", 6332=>X"0000003b0000003b0000003b0000003b", 6333=>X"0000003b0000003b0000003b0000003b", 6334=>X"0000003b0000003b0000003b0000003b", 
6335=>X"0000003b0000003b0000003b0000003b", 6336=>X"0000003b0000003b0000003b0000003b", 6337=>X"0000003b0000003b0000003b0000003b", 6338=>X"0000003b0000003b0000003b0000003b", 6339=>X"0000003b0000003b0000003b0000003b", 
6340=>X"0000003b0000003b0000003b0000003b", 6341=>X"0000003b0000003b0000003b0000003b", 6342=>X"0000003b0000003b0000003b0000003b", 6343=>X"0000003b0000003b0000003b0000003b", 6344=>X"0000003b0000003b0000003b0000003b", 
6345=>X"0000003b0000003b0000003b0000003b", 6346=>X"0000003b0000003b0000003b0000003b", 6347=>X"0000003b0000003b0000003b0000003b", 6348=>X"0000003b0000003b0000003b0000003b", 6349=>X"0000003b0000003b0000003b0000003b", 
6350=>X"0000003b0000003b0000003b0000003b", 6351=>X"0000003a0000003a0000003a0000003a", 6352=>X"0000003a0000003a0000003a0000003a", 6353=>X"0000003a0000003a0000003a0000003a", 6354=>X"0000003a0000003a0000003a0000003a", 
6355=>X"0000003a0000003a0000003a0000003a", 6356=>X"0000003a0000003a0000003a0000003a", 6357=>X"0000003a0000003a0000003a0000003a", 6358=>X"0000003a0000003a0000003a0000003a", 6359=>X"0000003a0000003a0000003a0000003a", 
6360=>X"0000003a0000003a0000003a0000003a", 6361=>X"0000003a0000003a0000003a0000003a", 6362=>X"0000003a0000003a0000003a0000003a", 6363=>X"0000003a0000003a0000003a0000003a", 6364=>X"0000003a0000003a0000003a0000003a", 
6365=>X"0000003a0000003a0000003a0000003a", 6366=>X"0000003a0000003a0000003a0000003a", 6367=>X"0000003a0000003a0000003a0000003a", 6368=>X"0000003a0000003a0000003a0000003a", 6369=>X"0000003a0000003a0000003a0000003a", 
6370=>X"0000003a0000003a0000003a0000003a", 6371=>X"0000003a0000003a0000003a0000003a", 6372=>X"0000003a0000003a0000003a0000003a", 6373=>X"0000003a0000003a0000003a0000003a", 6374=>X"0000003a0000003a0000003a0000003a", 
6375=>X"0000003a0000003a0000003a0000003a", 6376=>X"0000003a0000003a0000003a0000003a", 6377=>X"0000003a0000003a0000003a0000003a", 6378=>X"0000003a0000003a0000003a0000003a", 6379=>X"0000003a0000003a0000003a0000003a", 
6380=>X"0000003a0000003a0000003a0000003a", 6381=>X"0000003a0000003a0000003a0000003a", 6382=>X"0000003a0000003a0000003a0000003a", 6383=>X"0000003a0000003a0000003a0000003a", 6384=>X"0000003a0000003a0000003a0000003a", 
6385=>X"0000003a0000003a0000003a0000003a", 6386=>X"0000003a0000003a0000003a0000003a", 6387=>X"0000003a0000003a0000003a0000003a", 6388=>X"0000003a0000003a0000003a0000003a", 6389=>X"0000003a0000003a0000003a0000003a", 
6390=>X"0000003a0000003a0000003a0000003a", 6391=>X"0000003a0000003a0000003a0000003a", 6392=>X"0000003a0000003a0000003a0000003a", 6393=>X"0000003a0000003a0000003a0000003a", 6394=>X"0000003a0000003a0000003a0000003a", 
6395=>X"0000003a0000003a0000003a0000003a", 6396=>X"0000003a0000003a0000003a0000003a", 6397=>X"0000003a0000003a0000003a0000003a", 6398=>X"0000003a0000003a0000003a0000003a", 6399=>X"0000003a0000003a0000003a0000003a", 
6400=>X"0000003a0000003a0000003a0000003a", 6401=>X"0000003a0000003a0000003a0000003a", 6402=>X"0000003a0000003a0000003a0000003a", 6403=>X"0000003a0000003a0000003a0000003a", 6404=>X"0000003a0000003a0000003a0000003a", 
6405=>X"0000003a0000003a0000003a0000003a", 6406=>X"0000003a0000003a0000003a0000003a", 6407=>X"0000003a0000003a0000003a0000003a", 6408=>X"0000003a0000003a0000003a0000003a", 6409=>X"0000003a0000003a0000003a0000003a", 
6410=>X"0000003a0000003a0000003a0000003a", 6411=>X"0000003a0000003a0000003a0000003a", 6412=>X"0000003a0000003a0000003a0000003a", 6413=>X"0000003a0000003a0000003a0000003a", 6414=>X"0000003a0000003a0000003a0000003a", 
6415=>X"0000003a0000003a0000003a0000003a", 6416=>X"0000003a0000003a0000003a0000003a", 6417=>X"0000003a0000003a0000003a0000003a", 6418=>X"0000003a0000003a0000003a0000003a", 6419=>X"0000003a0000003a0000003a0000003a", 
6420=>X"0000003a0000003a0000003a0000003a", 6421=>X"0000003a0000003a0000003a0000003a", 6422=>X"0000003a0000003a0000003a0000003a", 6423=>X"0000003a0000003a0000003a0000003a", 6424=>X"0000003a0000003a0000003a0000003a", 
6425=>X"0000003a0000003a0000003a0000003a", 6426=>X"0000003a0000003a0000003a0000003a", 6427=>X"0000003a0000003a0000003a0000003a", 6428=>X"0000003a0000003a0000003a0000003a", 6429=>X"00000039000000390000003900000039", 
6430=>X"00000039000000390000003900000039", 6431=>X"00000039000000390000003900000039", 6432=>X"00000039000000390000003900000039", 6433=>X"00000039000000390000003900000039", 6434=>X"00000039000000390000003900000039", 
6435=>X"00000039000000390000003900000039", 6436=>X"00000039000000390000003900000039", 6437=>X"00000039000000390000003900000039", 6438=>X"00000039000000390000003900000039", 6439=>X"00000039000000390000003900000039", 
6440=>X"00000039000000390000003900000039", 6441=>X"00000039000000390000003900000039", 6442=>X"00000039000000390000003900000039", 6443=>X"00000039000000390000003900000039", 6444=>X"00000039000000390000003900000039", 
6445=>X"00000039000000390000003900000039", 6446=>X"00000039000000390000003900000039", 6447=>X"00000039000000390000003900000039", 6448=>X"00000039000000390000003900000039", 6449=>X"00000039000000390000003900000039", 
6450=>X"00000039000000390000003900000039", 6451=>X"00000039000000390000003900000039", 6452=>X"00000039000000390000003900000039", 6453=>X"00000039000000390000003900000039", 6454=>X"00000039000000390000003900000039", 
6455=>X"00000039000000390000003900000039", 6456=>X"00000039000000390000003900000039", 6457=>X"00000039000000390000003900000039", 6458=>X"00000039000000390000003900000039", 6459=>X"00000039000000390000003900000039", 
6460=>X"00000039000000390000003900000039", 6461=>X"00000039000000390000003900000039", 6462=>X"00000039000000390000003900000039", 6463=>X"00000039000000390000003900000039", 6464=>X"00000039000000390000003900000039", 
6465=>X"00000039000000390000003900000039", 6466=>X"00000039000000390000003900000039", 6467=>X"00000039000000390000003900000039", 6468=>X"00000039000000390000003900000039", 6469=>X"00000039000000390000003900000039", 
6470=>X"00000039000000390000003900000039", 6471=>X"00000039000000390000003900000039", 6472=>X"00000039000000390000003900000039", 6473=>X"00000039000000390000003900000039", 6474=>X"00000039000000390000003900000039", 
6475=>X"00000039000000390000003900000039", 6476=>X"00000039000000390000003900000039", 6477=>X"00000039000000390000003900000039", 6478=>X"00000039000000390000003900000039", 6479=>X"00000039000000390000003900000039", 
6480=>X"00000039000000390000003900000039", 6481=>X"00000039000000390000003900000039", 6482=>X"00000039000000390000003900000039", 6483=>X"00000039000000390000003900000039", 6484=>X"00000039000000390000003900000039", 
6485=>X"00000039000000390000003900000039", 6486=>X"00000039000000390000003900000039", 6487=>X"00000039000000390000003900000039", 6488=>X"00000039000000390000003900000039", 6489=>X"00000039000000390000003900000039", 
6490=>X"00000039000000390000003900000039", 6491=>X"00000039000000390000003900000039", 6492=>X"00000039000000390000003900000039", 6493=>X"00000039000000390000003900000039", 6494=>X"00000039000000390000003900000039", 
6495=>X"00000039000000390000003900000039", 6496=>X"00000039000000390000003900000039", 6497=>X"00000039000000390000003900000039", 6498=>X"00000039000000390000003900000039", 6499=>X"00000039000000390000003900000039", 
6500=>X"00000039000000390000003900000039", 6501=>X"00000039000000390000003900000039", 6502=>X"00000039000000390000003900000039", 6503=>X"00000039000000390000003900000039", 6504=>X"00000039000000390000003900000039", 
6505=>X"00000039000000390000003900000039", 6506=>X"00000039000000390000003900000039", 6507=>X"00000039000000390000003900000039", 6508=>X"00000039000000390000003900000039", 6509=>X"00000038000000380000003900000039", 
6510=>X"00000038000000380000003800000038", 6511=>X"00000038000000380000003800000038", 6512=>X"00000038000000380000003800000038", 6513=>X"00000038000000380000003800000038", 6514=>X"00000038000000380000003800000038", 
6515=>X"00000038000000380000003800000038", 6516=>X"00000038000000380000003800000038", 6517=>X"00000038000000380000003800000038", 6518=>X"00000038000000380000003800000038", 6519=>X"00000038000000380000003800000038", 
6520=>X"00000038000000380000003800000038", 6521=>X"00000038000000380000003800000038", 6522=>X"00000038000000380000003800000038", 6523=>X"00000038000000380000003800000038", 6524=>X"00000038000000380000003800000038", 
6525=>X"00000038000000380000003800000038", 6526=>X"00000038000000380000003800000038", 6527=>X"00000038000000380000003800000038", 6528=>X"00000038000000380000003800000038", 6529=>X"00000038000000380000003800000038", 
6530=>X"00000038000000380000003800000038", 6531=>X"00000038000000380000003800000038", 6532=>X"00000038000000380000003800000038", 6533=>X"00000038000000380000003800000038", 6534=>X"00000038000000380000003800000038", 
6535=>X"00000038000000380000003800000038", 6536=>X"00000038000000380000003800000038", 6537=>X"00000038000000380000003800000038", 6538=>X"00000038000000380000003800000038", 6539=>X"00000038000000380000003800000038", 
6540=>X"00000038000000380000003800000038", 6541=>X"00000038000000380000003800000038", 6542=>X"00000038000000380000003800000038", 6543=>X"00000038000000380000003800000038", 6544=>X"00000038000000380000003800000038", 
6545=>X"00000038000000380000003800000038", 6546=>X"00000038000000380000003800000038", 6547=>X"00000038000000380000003800000038", 6548=>X"00000038000000380000003800000038", 6549=>X"00000038000000380000003800000038", 
6550=>X"00000038000000380000003800000038", 6551=>X"00000038000000380000003800000038", 6552=>X"00000038000000380000003800000038", 6553=>X"00000038000000380000003800000038", 6554=>X"00000038000000380000003800000038", 
6555=>X"00000038000000380000003800000038", 6556=>X"00000038000000380000003800000038", 6557=>X"00000038000000380000003800000038", 6558=>X"00000038000000380000003800000038", 6559=>X"00000038000000380000003800000038", 
6560=>X"00000038000000380000003800000038", 6561=>X"00000038000000380000003800000038", 6562=>X"00000038000000380000003800000038", 6563=>X"00000038000000380000003800000038", 6564=>X"00000038000000380000003800000038", 
6565=>X"00000038000000380000003800000038", 6566=>X"00000038000000380000003800000038", 6567=>X"00000038000000380000003800000038", 6568=>X"00000038000000380000003800000038", 6569=>X"00000038000000380000003800000038", 
6570=>X"00000038000000380000003800000038", 6571=>X"00000038000000380000003800000038", 6572=>X"00000038000000380000003800000038", 6573=>X"00000038000000380000003800000038", 6574=>X"00000038000000380000003800000038", 
6575=>X"00000038000000380000003800000038", 6576=>X"00000038000000380000003800000038", 6577=>X"00000038000000380000003800000038", 6578=>X"00000038000000380000003800000038", 6579=>X"00000038000000380000003800000038", 
6580=>X"00000038000000380000003800000038", 6581=>X"00000038000000380000003800000038", 6582=>X"00000038000000380000003800000038", 6583=>X"00000038000000380000003800000038", 6584=>X"00000038000000380000003800000038", 
6585=>X"00000038000000380000003800000038", 6586=>X"00000038000000380000003800000038", 6587=>X"00000038000000380000003800000038", 6588=>X"00000038000000380000003800000038", 6589=>X"00000038000000380000003800000038", 
6590=>X"00000038000000380000003800000038", 6591=>X"00000038000000380000003800000038", 6592=>X"00000038000000380000003800000038", 6593=>X"00000037000000370000003700000038", 6594=>X"00000037000000370000003700000037", 
6595=>X"00000037000000370000003700000037", 6596=>X"00000037000000370000003700000037", 6597=>X"00000037000000370000003700000037", 6598=>X"00000037000000370000003700000037", 6599=>X"00000037000000370000003700000037", 
6600=>X"00000037000000370000003700000037", 6601=>X"00000037000000370000003700000037", 6602=>X"00000037000000370000003700000037", 6603=>X"00000037000000370000003700000037", 6604=>X"00000037000000370000003700000037", 
6605=>X"00000037000000370000003700000037", 6606=>X"00000037000000370000003700000037", 6607=>X"00000037000000370000003700000037", 6608=>X"00000037000000370000003700000037", 6609=>X"00000037000000370000003700000037", 
6610=>X"00000037000000370000003700000037", 6611=>X"00000037000000370000003700000037", 6612=>X"00000037000000370000003700000037", 6613=>X"00000037000000370000003700000037", 6614=>X"00000037000000370000003700000037", 
6615=>X"00000037000000370000003700000037", 6616=>X"00000037000000370000003700000037", 6617=>X"00000037000000370000003700000037", 6618=>X"00000037000000370000003700000037", 6619=>X"00000037000000370000003700000037", 
6620=>X"00000037000000370000003700000037", 6621=>X"00000037000000370000003700000037", 6622=>X"00000037000000370000003700000037", 6623=>X"00000037000000370000003700000037", 6624=>X"00000037000000370000003700000037", 
6625=>X"00000037000000370000003700000037", 6626=>X"00000037000000370000003700000037", 6627=>X"00000037000000370000003700000037", 6628=>X"00000037000000370000003700000037", 6629=>X"00000037000000370000003700000037", 
6630=>X"00000037000000370000003700000037", 6631=>X"00000037000000370000003700000037", 6632=>X"00000037000000370000003700000037", 6633=>X"00000037000000370000003700000037", 6634=>X"00000037000000370000003700000037", 
6635=>X"00000037000000370000003700000037", 6636=>X"00000037000000370000003700000037", 6637=>X"00000037000000370000003700000037", 6638=>X"00000037000000370000003700000037", 6639=>X"00000037000000370000003700000037", 
6640=>X"00000037000000370000003700000037", 6641=>X"00000037000000370000003700000037", 6642=>X"00000037000000370000003700000037", 6643=>X"00000037000000370000003700000037", 6644=>X"00000037000000370000003700000037", 
6645=>X"00000037000000370000003700000037", 6646=>X"00000037000000370000003700000037", 6647=>X"00000037000000370000003700000037", 6648=>X"00000037000000370000003700000037", 6649=>X"00000037000000370000003700000037", 
6650=>X"00000037000000370000003700000037", 6651=>X"00000037000000370000003700000037", 6652=>X"00000037000000370000003700000037", 6653=>X"00000037000000370000003700000037", 6654=>X"00000037000000370000003700000037", 
6655=>X"00000037000000370000003700000037", 6656=>X"00000037000000370000003700000037", 6657=>X"00000037000000370000003700000037", 6658=>X"00000037000000370000003700000037", 6659=>X"00000037000000370000003700000037", 
6660=>X"00000037000000370000003700000037", 6661=>X"00000037000000370000003700000037", 6662=>X"00000037000000370000003700000037", 6663=>X"00000037000000370000003700000037", 6664=>X"00000037000000370000003700000037", 
6665=>X"00000037000000370000003700000037", 6666=>X"00000037000000370000003700000037", 6667=>X"00000037000000370000003700000037", 6668=>X"00000037000000370000003700000037", 6669=>X"00000037000000370000003700000037", 
6670=>X"00000037000000370000003700000037", 6671=>X"00000037000000370000003700000037", 6672=>X"00000037000000370000003700000037", 6673=>X"00000037000000370000003700000037", 6674=>X"00000037000000370000003700000037", 
6675=>X"00000037000000370000003700000037", 6676=>X"00000037000000370000003700000037", 6677=>X"00000037000000370000003700000037", 6678=>X"00000037000000370000003700000037", 6679=>X"00000036000000370000003700000037", 
6680=>X"00000036000000360000003600000036", 6681=>X"00000036000000360000003600000036", 6682=>X"00000036000000360000003600000036", 6683=>X"00000036000000360000003600000036", 6684=>X"00000036000000360000003600000036", 
6685=>X"00000036000000360000003600000036", 6686=>X"00000036000000360000003600000036", 6687=>X"00000036000000360000003600000036", 6688=>X"00000036000000360000003600000036", 6689=>X"00000036000000360000003600000036", 
6690=>X"00000036000000360000003600000036", 6691=>X"00000036000000360000003600000036", 6692=>X"00000036000000360000003600000036", 6693=>X"00000036000000360000003600000036", 6694=>X"00000036000000360000003600000036", 
6695=>X"00000036000000360000003600000036", 6696=>X"00000036000000360000003600000036", 6697=>X"00000036000000360000003600000036", 6698=>X"00000036000000360000003600000036", 6699=>X"00000036000000360000003600000036", 
6700=>X"00000036000000360000003600000036", 6701=>X"00000036000000360000003600000036", 6702=>X"00000036000000360000003600000036", 6703=>X"00000036000000360000003600000036", 6704=>X"00000036000000360000003600000036", 
6705=>X"00000036000000360000003600000036", 6706=>X"00000036000000360000003600000036", 6707=>X"00000036000000360000003600000036", 6708=>X"00000036000000360000003600000036", 6709=>X"00000036000000360000003600000036", 
6710=>X"00000036000000360000003600000036", 6711=>X"00000036000000360000003600000036", 6712=>X"00000036000000360000003600000036", 6713=>X"00000036000000360000003600000036", 6714=>X"00000036000000360000003600000036", 
6715=>X"00000036000000360000003600000036", 6716=>X"00000036000000360000003600000036", 6717=>X"00000036000000360000003600000036", 6718=>X"00000036000000360000003600000036", 6719=>X"00000036000000360000003600000036", 
6720=>X"00000036000000360000003600000036", 6721=>X"00000036000000360000003600000036", 6722=>X"00000036000000360000003600000036", 6723=>X"00000036000000360000003600000036", 6724=>X"00000036000000360000003600000036", 
6725=>X"00000036000000360000003600000036", 6726=>X"00000036000000360000003600000036", 6727=>X"00000036000000360000003600000036", 6728=>X"00000036000000360000003600000036", 6729=>X"00000036000000360000003600000036", 
6730=>X"00000036000000360000003600000036", 6731=>X"00000036000000360000003600000036", 6732=>X"00000036000000360000003600000036", 6733=>X"00000036000000360000003600000036", 6734=>X"00000036000000360000003600000036", 
6735=>X"00000036000000360000003600000036", 6736=>X"00000036000000360000003600000036", 6737=>X"00000036000000360000003600000036", 6738=>X"00000036000000360000003600000036", 6739=>X"00000036000000360000003600000036", 
6740=>X"00000036000000360000003600000036", 6741=>X"00000036000000360000003600000036", 6742=>X"00000036000000360000003600000036", 6743=>X"00000036000000360000003600000036", 6744=>X"00000036000000360000003600000036", 
6745=>X"00000036000000360000003600000036", 6746=>X"00000036000000360000003600000036", 6747=>X"00000036000000360000003600000036", 6748=>X"00000036000000360000003600000036", 6749=>X"00000036000000360000003600000036", 
6750=>X"00000036000000360000003600000036", 6751=>X"00000036000000360000003600000036", 6752=>X"00000036000000360000003600000036", 6753=>X"00000036000000360000003600000036", 6754=>X"00000036000000360000003600000036", 
6755=>X"00000036000000360000003600000036", 6756=>X"00000036000000360000003600000036", 6757=>X"00000036000000360000003600000036", 6758=>X"00000036000000360000003600000036", 6759=>X"00000036000000360000003600000036", 
6760=>X"00000036000000360000003600000036", 6761=>X"00000036000000360000003600000036", 6762=>X"00000036000000360000003600000036", 6763=>X"00000036000000360000003600000036", 6764=>X"00000036000000360000003600000036", 
6765=>X"00000036000000360000003600000036", 6766=>X"00000036000000360000003600000036", 6767=>X"00000036000000360000003600000036", 6768=>X"00000036000000360000003600000036", 6769=>X"00000035000000360000003600000036", 
6770=>X"00000035000000350000003500000035", 6771=>X"00000035000000350000003500000035", 6772=>X"00000035000000350000003500000035", 6773=>X"00000035000000350000003500000035", 6774=>X"00000035000000350000003500000035", 
6775=>X"00000035000000350000003500000035", 6776=>X"00000035000000350000003500000035", 6777=>X"00000035000000350000003500000035", 6778=>X"00000035000000350000003500000035", 6779=>X"00000035000000350000003500000035", 
6780=>X"00000035000000350000003500000035", 6781=>X"00000035000000350000003500000035", 6782=>X"00000035000000350000003500000035", 6783=>X"00000035000000350000003500000035", 6784=>X"00000035000000350000003500000035", 
6785=>X"00000035000000350000003500000035", 6786=>X"00000035000000350000003500000035", 6787=>X"00000035000000350000003500000035", 6788=>X"00000035000000350000003500000035", 6789=>X"00000035000000350000003500000035", 
6790=>X"00000035000000350000003500000035", 6791=>X"00000035000000350000003500000035", 6792=>X"00000035000000350000003500000035", 6793=>X"00000035000000350000003500000035", 6794=>X"00000035000000350000003500000035", 
6795=>X"00000035000000350000003500000035", 6796=>X"00000035000000350000003500000035", 6797=>X"00000035000000350000003500000035", 6798=>X"00000035000000350000003500000035", 6799=>X"00000035000000350000003500000035", 
6800=>X"00000035000000350000003500000035", 6801=>X"00000035000000350000003500000035", 6802=>X"00000035000000350000003500000035", 6803=>X"00000035000000350000003500000035", 6804=>X"00000035000000350000003500000035", 
6805=>X"00000035000000350000003500000035", 6806=>X"00000035000000350000003500000035", 6807=>X"00000035000000350000003500000035", 6808=>X"00000035000000350000003500000035", 6809=>X"00000035000000350000003500000035", 
6810=>X"00000035000000350000003500000035", 6811=>X"00000035000000350000003500000035", 6812=>X"00000035000000350000003500000035", 6813=>X"00000035000000350000003500000035", 6814=>X"00000035000000350000003500000035", 
6815=>X"00000035000000350000003500000035", 6816=>X"00000035000000350000003500000035", 6817=>X"00000035000000350000003500000035", 6818=>X"00000035000000350000003500000035", 6819=>X"00000035000000350000003500000035", 
6820=>X"00000035000000350000003500000035", 6821=>X"00000035000000350000003500000035", 6822=>X"00000035000000350000003500000035", 6823=>X"00000035000000350000003500000035", 6824=>X"00000035000000350000003500000035", 
6825=>X"00000035000000350000003500000035", 6826=>X"00000035000000350000003500000035", 6827=>X"00000035000000350000003500000035", 6828=>X"00000035000000350000003500000035", 6829=>X"00000035000000350000003500000035", 
6830=>X"00000035000000350000003500000035", 6831=>X"00000035000000350000003500000035", 6832=>X"00000035000000350000003500000035", 6833=>X"00000035000000350000003500000035", 6834=>X"00000035000000350000003500000035", 
6835=>X"00000035000000350000003500000035", 6836=>X"00000035000000350000003500000035", 6837=>X"00000035000000350000003500000035", 6838=>X"00000035000000350000003500000035", 6839=>X"00000035000000350000003500000035", 
6840=>X"00000035000000350000003500000035", 6841=>X"00000035000000350000003500000035", 6842=>X"00000035000000350000003500000035", 6843=>X"00000035000000350000003500000035", 6844=>X"00000035000000350000003500000035", 
6845=>X"00000035000000350000003500000035", 6846=>X"00000035000000350000003500000035", 6847=>X"00000035000000350000003500000035", 6848=>X"00000035000000350000003500000035", 6849=>X"00000035000000350000003500000035", 
6850=>X"00000035000000350000003500000035", 6851=>X"00000035000000350000003500000035", 6852=>X"00000035000000350000003500000035", 6853=>X"00000035000000350000003500000035", 6854=>X"00000035000000350000003500000035", 
6855=>X"00000035000000350000003500000035", 6856=>X"00000035000000350000003500000035", 6857=>X"00000035000000350000003500000035", 6858=>X"00000035000000350000003500000035", 6859=>X"00000035000000350000003500000035", 
6860=>X"00000035000000350000003500000035", 6861=>X"00000035000000350000003500000035", 6862=>X"00000035000000350000003500000035", 6863=>X"00000034000000340000003400000034", 6864=>X"00000034000000340000003400000034", 
6865=>X"00000034000000340000003400000034", 6866=>X"00000034000000340000003400000034", 6867=>X"00000034000000340000003400000034", 6868=>X"00000034000000340000003400000034", 6869=>X"00000034000000340000003400000034", 
6870=>X"00000034000000340000003400000034", 6871=>X"00000034000000340000003400000034", 6872=>X"00000034000000340000003400000034", 6873=>X"00000034000000340000003400000034", 6874=>X"00000034000000340000003400000034", 
6875=>X"00000034000000340000003400000034", 6876=>X"00000034000000340000003400000034", 6877=>X"00000034000000340000003400000034", 6878=>X"00000034000000340000003400000034", 6879=>X"00000034000000340000003400000034", 
6880=>X"00000034000000340000003400000034", 6881=>X"00000034000000340000003400000034", 6882=>X"00000034000000340000003400000034", 6883=>X"00000034000000340000003400000034", 6884=>X"00000034000000340000003400000034", 
6885=>X"00000034000000340000003400000034", 6886=>X"00000034000000340000003400000034", 6887=>X"00000034000000340000003400000034", 6888=>X"00000034000000340000003400000034", 6889=>X"00000034000000340000003400000034", 
6890=>X"00000034000000340000003400000034", 6891=>X"00000034000000340000003400000034", 6892=>X"00000034000000340000003400000034", 6893=>X"00000034000000340000003400000034", 6894=>X"00000034000000340000003400000034", 
6895=>X"00000034000000340000003400000034", 6896=>X"00000034000000340000003400000034", 6897=>X"00000034000000340000003400000034", 6898=>X"00000034000000340000003400000034", 6899=>X"00000034000000340000003400000034", 
6900=>X"00000034000000340000003400000034", 6901=>X"00000034000000340000003400000034", 6902=>X"00000034000000340000003400000034", 6903=>X"00000034000000340000003400000034", 6904=>X"00000034000000340000003400000034", 
6905=>X"00000034000000340000003400000034", 6906=>X"00000034000000340000003400000034", 6907=>X"00000034000000340000003400000034", 6908=>X"00000034000000340000003400000034", 6909=>X"00000034000000340000003400000034", 
6910=>X"00000034000000340000003400000034", 6911=>X"00000034000000340000003400000034", 6912=>X"00000034000000340000003400000034", 6913=>X"00000034000000340000003400000034", 6914=>X"00000034000000340000003400000034", 
6915=>X"00000034000000340000003400000034", 6916=>X"00000034000000340000003400000034", 6917=>X"00000034000000340000003400000034", 6918=>X"00000034000000340000003400000034", 6919=>X"00000034000000340000003400000034", 
6920=>X"00000034000000340000003400000034", 6921=>X"00000034000000340000003400000034", 6922=>X"00000034000000340000003400000034", 6923=>X"00000034000000340000003400000034", 6924=>X"00000034000000340000003400000034", 
6925=>X"00000034000000340000003400000034", 6926=>X"00000034000000340000003400000034", 6927=>X"00000034000000340000003400000034", 6928=>X"00000034000000340000003400000034", 6929=>X"00000034000000340000003400000034", 
6930=>X"00000034000000340000003400000034", 6931=>X"00000034000000340000003400000034", 6932=>X"00000034000000340000003400000034", 6933=>X"00000034000000340000003400000034", 6934=>X"00000034000000340000003400000034", 
6935=>X"00000034000000340000003400000034", 6936=>X"00000034000000340000003400000034", 6937=>X"00000034000000340000003400000034", 6938=>X"00000034000000340000003400000034", 6939=>X"00000034000000340000003400000034", 
6940=>X"00000034000000340000003400000034", 6941=>X"00000034000000340000003400000034", 6942=>X"00000034000000340000003400000034", 6943=>X"00000034000000340000003400000034", 6944=>X"00000034000000340000003400000034", 
6945=>X"00000034000000340000003400000034", 6946=>X"00000034000000340000003400000034", 6947=>X"00000034000000340000003400000034", 6948=>X"00000034000000340000003400000034", 6949=>X"00000034000000340000003400000034", 
6950=>X"00000034000000340000003400000034", 6951=>X"00000034000000340000003400000034", 6952=>X"00000034000000340000003400000034", 6953=>X"00000034000000340000003400000034", 6954=>X"00000034000000340000003400000034", 
6955=>X"00000034000000340000003400000034", 6956=>X"00000034000000340000003400000034", 6957=>X"00000034000000340000003400000034", 6958=>X"00000034000000340000003400000034", 6959=>X"00000034000000340000003400000034", 
6960=>X"00000033000000330000003300000033", 6961=>X"00000033000000330000003300000033", 6962=>X"00000033000000330000003300000033", 6963=>X"00000033000000330000003300000033", 6964=>X"00000033000000330000003300000033", 
6965=>X"00000033000000330000003300000033", 6966=>X"00000033000000330000003300000033", 6967=>X"00000033000000330000003300000033", 6968=>X"00000033000000330000003300000033", 6969=>X"00000033000000330000003300000033", 
6970=>X"00000033000000330000003300000033", 6971=>X"00000033000000330000003300000033", 6972=>X"00000033000000330000003300000033", 6973=>X"00000033000000330000003300000033", 6974=>X"00000033000000330000003300000033", 
6975=>X"00000033000000330000003300000033", 6976=>X"00000033000000330000003300000033", 6977=>X"00000033000000330000003300000033", 6978=>X"00000033000000330000003300000033", 6979=>X"00000033000000330000003300000033", 
6980=>X"00000033000000330000003300000033", 6981=>X"00000033000000330000003300000033", 6982=>X"00000033000000330000003300000033", 6983=>X"00000033000000330000003300000033", 6984=>X"00000033000000330000003300000033", 
6985=>X"00000033000000330000003300000033", 6986=>X"00000033000000330000003300000033", 6987=>X"00000033000000330000003300000033", 6988=>X"00000033000000330000003300000033", 6989=>X"00000033000000330000003300000033", 
6990=>X"00000033000000330000003300000033", 6991=>X"00000033000000330000003300000033", 6992=>X"00000033000000330000003300000033", 6993=>X"00000033000000330000003300000033", 6994=>X"00000033000000330000003300000033", 
6995=>X"00000033000000330000003300000033", 6996=>X"00000033000000330000003300000033", 6997=>X"00000033000000330000003300000033", 6998=>X"00000033000000330000003300000033", 6999=>X"00000033000000330000003300000033", 
7000=>X"00000033000000330000003300000033", 7001=>X"00000033000000330000003300000033", 7002=>X"00000033000000330000003300000033", 7003=>X"00000033000000330000003300000033", 7004=>X"00000033000000330000003300000033", 
7005=>X"00000033000000330000003300000033", 7006=>X"00000033000000330000003300000033", 7007=>X"00000033000000330000003300000033", 7008=>X"00000033000000330000003300000033", 7009=>X"00000033000000330000003300000033", 
7010=>X"00000033000000330000003300000033", 7011=>X"00000033000000330000003300000033", 7012=>X"00000033000000330000003300000033", 7013=>X"00000033000000330000003300000033", 7014=>X"00000033000000330000003300000033", 
7015=>X"00000033000000330000003300000033", 7016=>X"00000033000000330000003300000033", 7017=>X"00000033000000330000003300000033", 7018=>X"00000033000000330000003300000033", 7019=>X"00000033000000330000003300000033", 
7020=>X"00000033000000330000003300000033", 7021=>X"00000033000000330000003300000033", 7022=>X"00000033000000330000003300000033", 7023=>X"00000033000000330000003300000033", 7024=>X"00000033000000330000003300000033", 
7025=>X"00000033000000330000003300000033", 7026=>X"00000033000000330000003300000033", 7027=>X"00000033000000330000003300000033", 7028=>X"00000033000000330000003300000033", 7029=>X"00000033000000330000003300000033", 
7030=>X"00000033000000330000003300000033", 7031=>X"00000033000000330000003300000033", 7032=>X"00000033000000330000003300000033", 7033=>X"00000033000000330000003300000033", 7034=>X"00000033000000330000003300000033", 
7035=>X"00000033000000330000003300000033", 7036=>X"00000033000000330000003300000033", 7037=>X"00000033000000330000003300000033", 7038=>X"00000033000000330000003300000033", 7039=>X"00000033000000330000003300000033", 
7040=>X"00000033000000330000003300000033", 7041=>X"00000033000000330000003300000033", 7042=>X"00000033000000330000003300000033", 7043=>X"00000033000000330000003300000033", 7044=>X"00000033000000330000003300000033", 
7045=>X"00000033000000330000003300000033", 7046=>X"00000033000000330000003300000033", 7047=>X"00000033000000330000003300000033", 7048=>X"00000033000000330000003300000033", 7049=>X"00000033000000330000003300000033", 
7050=>X"00000033000000330000003300000033", 7051=>X"00000033000000330000003300000033", 7052=>X"00000033000000330000003300000033", 7053=>X"00000033000000330000003300000033", 7054=>X"00000033000000330000003300000033", 
7055=>X"00000033000000330000003300000033", 7056=>X"00000033000000330000003300000033", 7057=>X"00000033000000330000003300000033", 7058=>X"00000033000000330000003300000033", 7059=>X"00000033000000330000003300000033", 
7060=>X"00000032000000330000003300000033", 7061=>X"00000032000000320000003200000032", 7062=>X"00000032000000320000003200000032", 7063=>X"00000032000000320000003200000032", 7064=>X"00000032000000320000003200000032", 
7065=>X"00000032000000320000003200000032", 7066=>X"00000032000000320000003200000032", 7067=>X"00000032000000320000003200000032", 7068=>X"00000032000000320000003200000032", 7069=>X"00000032000000320000003200000032", 
7070=>X"00000032000000320000003200000032", 7071=>X"00000032000000320000003200000032", 7072=>X"00000032000000320000003200000032", 7073=>X"00000032000000320000003200000032", 7074=>X"00000032000000320000003200000032", 
7075=>X"00000032000000320000003200000032", 7076=>X"00000032000000320000003200000032", 7077=>X"00000032000000320000003200000032", 7078=>X"00000032000000320000003200000032", 7079=>X"00000032000000320000003200000032", 
7080=>X"00000032000000320000003200000032", 7081=>X"00000032000000320000003200000032", 7082=>X"00000032000000320000003200000032", 7083=>X"00000032000000320000003200000032", 7084=>X"00000032000000320000003200000032", 
7085=>X"00000032000000320000003200000032", 7086=>X"00000032000000320000003200000032", 7087=>X"00000032000000320000003200000032", 7088=>X"00000032000000320000003200000032", 7089=>X"00000032000000320000003200000032", 
7090=>X"00000032000000320000003200000032", 7091=>X"00000032000000320000003200000032", 7092=>X"00000032000000320000003200000032", 7093=>X"00000032000000320000003200000032", 7094=>X"00000032000000320000003200000032", 
7095=>X"00000032000000320000003200000032", 7096=>X"00000032000000320000003200000032", 7097=>X"00000032000000320000003200000032", 7098=>X"00000032000000320000003200000032", 7099=>X"00000032000000320000003200000032", 
7100=>X"00000032000000320000003200000032", 7101=>X"00000032000000320000003200000032", 7102=>X"00000032000000320000003200000032", 7103=>X"00000032000000320000003200000032", 7104=>X"00000032000000320000003200000032", 
7105=>X"00000032000000320000003200000032", 7106=>X"00000032000000320000003200000032", 7107=>X"00000032000000320000003200000032", 7108=>X"00000032000000320000003200000032", 7109=>X"00000032000000320000003200000032", 
7110=>X"00000032000000320000003200000032", 7111=>X"00000032000000320000003200000032", 7112=>X"00000032000000320000003200000032", 7113=>X"00000032000000320000003200000032", 7114=>X"00000032000000320000003200000032", 
7115=>X"00000032000000320000003200000032", 7116=>X"00000032000000320000003200000032", 7117=>X"00000032000000320000003200000032", 7118=>X"00000032000000320000003200000032", 7119=>X"00000032000000320000003200000032", 
7120=>X"00000032000000320000003200000032", 7121=>X"00000032000000320000003200000032", 7122=>X"00000032000000320000003200000032", 7123=>X"00000032000000320000003200000032", 7124=>X"00000032000000320000003200000032", 
7125=>X"00000032000000320000003200000032", 7126=>X"00000032000000320000003200000032", 7127=>X"00000032000000320000003200000032", 7128=>X"00000032000000320000003200000032", 7129=>X"00000032000000320000003200000032", 
7130=>X"00000032000000320000003200000032", 7131=>X"00000032000000320000003200000032", 7132=>X"00000032000000320000003200000032", 7133=>X"00000032000000320000003200000032", 7134=>X"00000032000000320000003200000032", 
7135=>X"00000032000000320000003200000032", 7136=>X"00000032000000320000003200000032", 7137=>X"00000032000000320000003200000032", 7138=>X"00000032000000320000003200000032", 7139=>X"00000032000000320000003200000032", 
7140=>X"00000032000000320000003200000032", 7141=>X"00000032000000320000003200000032", 7142=>X"00000032000000320000003200000032", 7143=>X"00000032000000320000003200000032", 7144=>X"00000032000000320000003200000032", 
7145=>X"00000032000000320000003200000032", 7146=>X"00000032000000320000003200000032", 7147=>X"00000032000000320000003200000032", 7148=>X"00000032000000320000003200000032", 7149=>X"00000032000000320000003200000032", 
7150=>X"00000032000000320000003200000032", 7151=>X"00000032000000320000003200000032", 7152=>X"00000032000000320000003200000032", 7153=>X"00000032000000320000003200000032", 7154=>X"00000032000000320000003200000032", 
7155=>X"00000032000000320000003200000032", 7156=>X"00000032000000320000003200000032", 7157=>X"00000032000000320000003200000032", 7158=>X"00000032000000320000003200000032", 7159=>X"00000032000000320000003200000032", 
7160=>X"00000032000000320000003200000032", 7161=>X"00000032000000320000003200000032", 7162=>X"00000032000000320000003200000032", 7163=>X"00000032000000320000003200000032", 7164=>X"00000032000000320000003200000032", 
7165=>X"00000031000000320000003200000032", 7166=>X"00000031000000310000003100000031", 7167=>X"00000031000000310000003100000031", 7168=>X"00000031000000310000003100000031", 7169=>X"00000031000000310000003100000031", 
7170=>X"00000031000000310000003100000031", 7171=>X"00000031000000310000003100000031", 7172=>X"00000031000000310000003100000031", 7173=>X"00000031000000310000003100000031", 7174=>X"00000031000000310000003100000031", 
7175=>X"00000031000000310000003100000031", 7176=>X"00000031000000310000003100000031", 7177=>X"00000031000000310000003100000031", 7178=>X"00000031000000310000003100000031", 7179=>X"00000031000000310000003100000031", 
7180=>X"00000031000000310000003100000031", 7181=>X"00000031000000310000003100000031", 7182=>X"00000031000000310000003100000031", 7183=>X"00000031000000310000003100000031", 7184=>X"00000031000000310000003100000031", 
7185=>X"00000031000000310000003100000031", 7186=>X"00000031000000310000003100000031", 7187=>X"00000031000000310000003100000031", 7188=>X"00000031000000310000003100000031", 7189=>X"00000031000000310000003100000031", 
7190=>X"00000031000000310000003100000031", 7191=>X"00000031000000310000003100000031", 7192=>X"00000031000000310000003100000031", 7193=>X"00000031000000310000003100000031", 7194=>X"00000031000000310000003100000031", 
7195=>X"00000031000000310000003100000031", 7196=>X"00000031000000310000003100000031", 7197=>X"00000031000000310000003100000031", 7198=>X"00000031000000310000003100000031", 7199=>X"00000031000000310000003100000031", 
7200=>X"00000031000000310000003100000031", 7201=>X"00000031000000310000003100000031", 7202=>X"00000031000000310000003100000031", 7203=>X"00000031000000310000003100000031", 7204=>X"00000031000000310000003100000031", 
7205=>X"00000031000000310000003100000031", 7206=>X"00000031000000310000003100000031", 7207=>X"00000031000000310000003100000031", 7208=>X"00000031000000310000003100000031", 7209=>X"00000031000000310000003100000031", 
7210=>X"00000031000000310000003100000031", 7211=>X"00000031000000310000003100000031", 7212=>X"00000031000000310000003100000031", 7213=>X"00000031000000310000003100000031", 7214=>X"00000031000000310000003100000031", 
7215=>X"00000031000000310000003100000031", 7216=>X"00000031000000310000003100000031", 7217=>X"00000031000000310000003100000031", 7218=>X"00000031000000310000003100000031", 7219=>X"00000031000000310000003100000031", 
7220=>X"00000031000000310000003100000031", 7221=>X"00000031000000310000003100000031", 7222=>X"00000031000000310000003100000031", 7223=>X"00000031000000310000003100000031", 7224=>X"00000031000000310000003100000031", 
7225=>X"00000031000000310000003100000031", 7226=>X"00000031000000310000003100000031", 7227=>X"00000031000000310000003100000031", 7228=>X"00000031000000310000003100000031", 7229=>X"00000031000000310000003100000031", 
7230=>X"00000031000000310000003100000031", 7231=>X"00000031000000310000003100000031", 7232=>X"00000031000000310000003100000031", 7233=>X"00000031000000310000003100000031", 7234=>X"00000031000000310000003100000031", 
7235=>X"00000031000000310000003100000031", 7236=>X"00000031000000310000003100000031", 7237=>X"00000031000000310000003100000031", 7238=>X"00000031000000310000003100000031", 7239=>X"00000031000000310000003100000031", 
7240=>X"00000031000000310000003100000031", 7241=>X"00000031000000310000003100000031", 7242=>X"00000031000000310000003100000031", 7243=>X"00000031000000310000003100000031", 7244=>X"00000031000000310000003100000031", 
7245=>X"00000031000000310000003100000031", 7246=>X"00000031000000310000003100000031", 7247=>X"00000031000000310000003100000031", 7248=>X"00000031000000310000003100000031", 7249=>X"00000031000000310000003100000031", 
7250=>X"00000031000000310000003100000031", 7251=>X"00000031000000310000003100000031", 7252=>X"00000031000000310000003100000031", 7253=>X"00000031000000310000003100000031", 7254=>X"00000031000000310000003100000031", 
7255=>X"00000031000000310000003100000031", 7256=>X"00000031000000310000003100000031", 7257=>X"00000031000000310000003100000031", 7258=>X"00000031000000310000003100000031", 7259=>X"00000031000000310000003100000031", 
7260=>X"00000031000000310000003100000031", 7261=>X"00000031000000310000003100000031", 7262=>X"00000031000000310000003100000031", 7263=>X"00000031000000310000003100000031", 7264=>X"00000031000000310000003100000031", 
7265=>X"00000031000000310000003100000031", 7266=>X"00000031000000310000003100000031", 7267=>X"00000031000000310000003100000031", 7268=>X"00000031000000310000003100000031", 7269=>X"00000031000000310000003100000031", 
7270=>X"00000031000000310000003100000031", 7271=>X"00000031000000310000003100000031", 7272=>X"00000031000000310000003100000031", 7273=>X"00000031000000310000003100000031", 7274=>X"00000031000000310000003100000031", 
7275=>X"00000030000000300000003000000030", 7276=>X"00000030000000300000003000000030", 7277=>X"00000030000000300000003000000030", 7278=>X"00000030000000300000003000000030", 7279=>X"00000030000000300000003000000030", 
7280=>X"00000030000000300000003000000030", 7281=>X"00000030000000300000003000000030", 7282=>X"00000030000000300000003000000030", 7283=>X"00000030000000300000003000000030", 7284=>X"00000030000000300000003000000030", 
7285=>X"00000030000000300000003000000030", 7286=>X"00000030000000300000003000000030", 7287=>X"00000030000000300000003000000030", 7288=>X"00000030000000300000003000000030", 7289=>X"00000030000000300000003000000030", 
7290=>X"00000030000000300000003000000030", 7291=>X"00000030000000300000003000000030", 7292=>X"00000030000000300000003000000030", 7293=>X"00000030000000300000003000000030", 7294=>X"00000030000000300000003000000030", 
7295=>X"00000030000000300000003000000030", 7296=>X"00000030000000300000003000000030", 7297=>X"00000030000000300000003000000030", 7298=>X"00000030000000300000003000000030", 7299=>X"00000030000000300000003000000030", 
7300=>X"00000030000000300000003000000030", 7301=>X"00000030000000300000003000000030", 7302=>X"00000030000000300000003000000030", 7303=>X"00000030000000300000003000000030", 7304=>X"00000030000000300000003000000030", 
7305=>X"00000030000000300000003000000030", 7306=>X"00000030000000300000003000000030", 7307=>X"00000030000000300000003000000030", 7308=>X"00000030000000300000003000000030", 7309=>X"00000030000000300000003000000030", 
7310=>X"00000030000000300000003000000030", 7311=>X"00000030000000300000003000000030", 7312=>X"00000030000000300000003000000030", 7313=>X"00000030000000300000003000000030", 7314=>X"00000030000000300000003000000030", 
7315=>X"00000030000000300000003000000030", 7316=>X"00000030000000300000003000000030", 7317=>X"00000030000000300000003000000030", 7318=>X"00000030000000300000003000000030", 7319=>X"00000030000000300000003000000030", 
7320=>X"00000030000000300000003000000030", 7321=>X"00000030000000300000003000000030", 7322=>X"00000030000000300000003000000030", 7323=>X"00000030000000300000003000000030", 7324=>X"00000030000000300000003000000030", 
7325=>X"00000030000000300000003000000030", 7326=>X"00000030000000300000003000000030", 7327=>X"00000030000000300000003000000030", 7328=>X"00000030000000300000003000000030", 7329=>X"00000030000000300000003000000030", 
7330=>X"00000030000000300000003000000030", 7331=>X"00000030000000300000003000000030", 7332=>X"00000030000000300000003000000030", 7333=>X"00000030000000300000003000000030", 7334=>X"00000030000000300000003000000030", 
7335=>X"00000030000000300000003000000030", 7336=>X"00000030000000300000003000000030", 7337=>X"00000030000000300000003000000030", 7338=>X"00000030000000300000003000000030", 7339=>X"00000030000000300000003000000030", 
7340=>X"00000030000000300000003000000030", 7341=>X"00000030000000300000003000000030", 7342=>X"00000030000000300000003000000030", 7343=>X"00000030000000300000003000000030", 7344=>X"00000030000000300000003000000030", 
7345=>X"00000030000000300000003000000030", 7346=>X"00000030000000300000003000000030", 7347=>X"00000030000000300000003000000030", 7348=>X"00000030000000300000003000000030", 7349=>X"00000030000000300000003000000030", 
7350=>X"00000030000000300000003000000030", 7351=>X"00000030000000300000003000000030", 7352=>X"00000030000000300000003000000030", 7353=>X"00000030000000300000003000000030", 7354=>X"00000030000000300000003000000030", 
7355=>X"00000030000000300000003000000030", 7356=>X"00000030000000300000003000000030", 7357=>X"00000030000000300000003000000030", 7358=>X"00000030000000300000003000000030", 7359=>X"00000030000000300000003000000030", 
7360=>X"00000030000000300000003000000030", 7361=>X"00000030000000300000003000000030", 7362=>X"00000030000000300000003000000030", 7363=>X"00000030000000300000003000000030", 7364=>X"00000030000000300000003000000030", 
7365=>X"00000030000000300000003000000030", 7366=>X"00000030000000300000003000000030", 7367=>X"00000030000000300000003000000030", 7368=>X"00000030000000300000003000000030", 7369=>X"00000030000000300000003000000030", 
7370=>X"00000030000000300000003000000030", 7371=>X"00000030000000300000003000000030", 7372=>X"00000030000000300000003000000030", 7373=>X"00000030000000300000003000000030", 7374=>X"00000030000000300000003000000030", 
7375=>X"00000030000000300000003000000030", 7376=>X"00000030000000300000003000000030", 7377=>X"00000030000000300000003000000030", 7378=>X"00000030000000300000003000000030", 7379=>X"00000030000000300000003000000030", 
7380=>X"00000030000000300000003000000030", 7381=>X"00000030000000300000003000000030", 7382=>X"00000030000000300000003000000030", 7383=>X"00000030000000300000003000000030", 7384=>X"00000030000000300000003000000030", 
7385=>X"00000030000000300000003000000030", 7386=>X"00000030000000300000003000000030", 7387=>X"00000030000000300000003000000030", 7388=>X"0000002f000000300000003000000030", 7389=>X"0000002f0000002f0000002f0000002f", 
7390=>X"0000002f0000002f0000002f0000002f", 7391=>X"0000002f0000002f0000002f0000002f", 7392=>X"0000002f0000002f0000002f0000002f", 7393=>X"0000002f0000002f0000002f0000002f", 7394=>X"0000002f0000002f0000002f0000002f", 
7395=>X"0000002f0000002f0000002f0000002f", 7396=>X"0000002f0000002f0000002f0000002f", 7397=>X"0000002f0000002f0000002f0000002f", 7398=>X"0000002f0000002f0000002f0000002f", 7399=>X"0000002f0000002f0000002f0000002f", 
7400=>X"0000002f0000002f0000002f0000002f", 7401=>X"0000002f0000002f0000002f0000002f", 7402=>X"0000002f0000002f0000002f0000002f", 7403=>X"0000002f0000002f0000002f0000002f", 7404=>X"0000002f0000002f0000002f0000002f", 
7405=>X"0000002f0000002f0000002f0000002f", 7406=>X"0000002f0000002f0000002f0000002f", 7407=>X"0000002f0000002f0000002f0000002f", 7408=>X"0000002f0000002f0000002f0000002f", 7409=>X"0000002f0000002f0000002f0000002f", 
7410=>X"0000002f0000002f0000002f0000002f", 7411=>X"0000002f0000002f0000002f0000002f", 7412=>X"0000002f0000002f0000002f0000002f", 7413=>X"0000002f0000002f0000002f0000002f", 7414=>X"0000002f0000002f0000002f0000002f", 
7415=>X"0000002f0000002f0000002f0000002f", 7416=>X"0000002f0000002f0000002f0000002f", 7417=>X"0000002f0000002f0000002f0000002f", 7418=>X"0000002f0000002f0000002f0000002f", 7419=>X"0000002f0000002f0000002f0000002f", 
7420=>X"0000002f0000002f0000002f0000002f", 7421=>X"0000002f0000002f0000002f0000002f", 7422=>X"0000002f0000002f0000002f0000002f", 7423=>X"0000002f0000002f0000002f0000002f", 7424=>X"0000002f0000002f0000002f0000002f", 
7425=>X"0000002f0000002f0000002f0000002f", 7426=>X"0000002f0000002f0000002f0000002f", 7427=>X"0000002f0000002f0000002f0000002f", 7428=>X"0000002f0000002f0000002f0000002f", 7429=>X"0000002f0000002f0000002f0000002f", 
7430=>X"0000002f0000002f0000002f0000002f", 7431=>X"0000002f0000002f0000002f0000002f", 7432=>X"0000002f0000002f0000002f0000002f", 7433=>X"0000002f0000002f0000002f0000002f", 7434=>X"0000002f0000002f0000002f0000002f", 
7435=>X"0000002f0000002f0000002f0000002f", 7436=>X"0000002f0000002f0000002f0000002f", 7437=>X"0000002f0000002f0000002f0000002f", 7438=>X"0000002f0000002f0000002f0000002f", 7439=>X"0000002f0000002f0000002f0000002f", 
7440=>X"0000002f0000002f0000002f0000002f", 7441=>X"0000002f0000002f0000002f0000002f", 7442=>X"0000002f0000002f0000002f0000002f", 7443=>X"0000002f0000002f0000002f0000002f", 7444=>X"0000002f0000002f0000002f0000002f", 
7445=>X"0000002f0000002f0000002f0000002f", 7446=>X"0000002f0000002f0000002f0000002f", 7447=>X"0000002f0000002f0000002f0000002f", 7448=>X"0000002f0000002f0000002f0000002f", 7449=>X"0000002f0000002f0000002f0000002f", 
7450=>X"0000002f0000002f0000002f0000002f", 7451=>X"0000002f0000002f0000002f0000002f", 7452=>X"0000002f0000002f0000002f0000002f", 7453=>X"0000002f0000002f0000002f0000002f", 7454=>X"0000002f0000002f0000002f0000002f", 
7455=>X"0000002f0000002f0000002f0000002f", 7456=>X"0000002f0000002f0000002f0000002f", 7457=>X"0000002f0000002f0000002f0000002f", 7458=>X"0000002f0000002f0000002f0000002f", 7459=>X"0000002f0000002f0000002f0000002f", 
7460=>X"0000002f0000002f0000002f0000002f", 7461=>X"0000002f0000002f0000002f0000002f", 7462=>X"0000002f0000002f0000002f0000002f", 7463=>X"0000002f0000002f0000002f0000002f", 7464=>X"0000002f0000002f0000002f0000002f", 
7465=>X"0000002f0000002f0000002f0000002f", 7466=>X"0000002f0000002f0000002f0000002f", 7467=>X"0000002f0000002f0000002f0000002f", 7468=>X"0000002f0000002f0000002f0000002f", 7469=>X"0000002f0000002f0000002f0000002f", 
7470=>X"0000002f0000002f0000002f0000002f", 7471=>X"0000002f0000002f0000002f0000002f", 7472=>X"0000002f0000002f0000002f0000002f", 7473=>X"0000002f0000002f0000002f0000002f", 7474=>X"0000002f0000002f0000002f0000002f", 
7475=>X"0000002f0000002f0000002f0000002f", 7476=>X"0000002f0000002f0000002f0000002f", 7477=>X"0000002f0000002f0000002f0000002f", 7478=>X"0000002f0000002f0000002f0000002f", 7479=>X"0000002f0000002f0000002f0000002f", 
7480=>X"0000002f0000002f0000002f0000002f", 7481=>X"0000002f0000002f0000002f0000002f", 7482=>X"0000002f0000002f0000002f0000002f", 7483=>X"0000002f0000002f0000002f0000002f", 7484=>X"0000002f0000002f0000002f0000002f", 
7485=>X"0000002f0000002f0000002f0000002f", 7486=>X"0000002f0000002f0000002f0000002f", 7487=>X"0000002f0000002f0000002f0000002f", 7488=>X"0000002f0000002f0000002f0000002f", 7489=>X"0000002f0000002f0000002f0000002f", 
7490=>X"0000002f0000002f0000002f0000002f", 7491=>X"0000002f0000002f0000002f0000002f", 7492=>X"0000002f0000002f0000002f0000002f", 7493=>X"0000002f0000002f0000002f0000002f", 7494=>X"0000002f0000002f0000002f0000002f", 
7495=>X"0000002f0000002f0000002f0000002f", 7496=>X"0000002f0000002f0000002f0000002f", 7497=>X"0000002f0000002f0000002f0000002f", 7498=>X"0000002f0000002f0000002f0000002f", 7499=>X"0000002f0000002f0000002f0000002f", 
7500=>X"0000002f0000002f0000002f0000002f", 7501=>X"0000002f0000002f0000002f0000002f", 7502=>X"0000002f0000002f0000002f0000002f", 7503=>X"0000002f0000002f0000002f0000002f", 7504=>X"0000002f0000002f0000002f0000002f", 
7505=>X"0000002f0000002f0000002f0000002f", 7506=>X"0000002f0000002f0000002f0000002f", 7507=>X"0000002e0000002e0000002f0000002f", 7508=>X"0000002e0000002e0000002e0000002e", 7509=>X"0000002e0000002e0000002e0000002e", 
7510=>X"0000002e0000002e0000002e0000002e", 7511=>X"0000002e0000002e0000002e0000002e", 7512=>X"0000002e0000002e0000002e0000002e", 7513=>X"0000002e0000002e0000002e0000002e", 7514=>X"0000002e0000002e0000002e0000002e", 
7515=>X"0000002e0000002e0000002e0000002e", 7516=>X"0000002e0000002e0000002e0000002e", 7517=>X"0000002e0000002e0000002e0000002e", 7518=>X"0000002e0000002e0000002e0000002e", 7519=>X"0000002e0000002e0000002e0000002e", 
7520=>X"0000002e0000002e0000002e0000002e", 7521=>X"0000002e0000002e0000002e0000002e", 7522=>X"0000002e0000002e0000002e0000002e", 7523=>X"0000002e0000002e0000002e0000002e", 7524=>X"0000002e0000002e0000002e0000002e", 
7525=>X"0000002e0000002e0000002e0000002e", 7526=>X"0000002e0000002e0000002e0000002e", 7527=>X"0000002e0000002e0000002e0000002e", 7528=>X"0000002e0000002e0000002e0000002e", 7529=>X"0000002e0000002e0000002e0000002e", 
7530=>X"0000002e0000002e0000002e0000002e", 7531=>X"0000002e0000002e0000002e0000002e", 7532=>X"0000002e0000002e0000002e0000002e", 7533=>X"0000002e0000002e0000002e0000002e", 7534=>X"0000002e0000002e0000002e0000002e", 
7535=>X"0000002e0000002e0000002e0000002e", 7536=>X"0000002e0000002e0000002e0000002e", 7537=>X"0000002e0000002e0000002e0000002e", 7538=>X"0000002e0000002e0000002e0000002e", 7539=>X"0000002e0000002e0000002e0000002e", 
7540=>X"0000002e0000002e0000002e0000002e", 7541=>X"0000002e0000002e0000002e0000002e", 7542=>X"0000002e0000002e0000002e0000002e", 7543=>X"0000002e0000002e0000002e0000002e", 7544=>X"0000002e0000002e0000002e0000002e", 
7545=>X"0000002e0000002e0000002e0000002e", 7546=>X"0000002e0000002e0000002e0000002e", 7547=>X"0000002e0000002e0000002e0000002e", 7548=>X"0000002e0000002e0000002e0000002e", 7549=>X"0000002e0000002e0000002e0000002e", 
7550=>X"0000002e0000002e0000002e0000002e", 7551=>X"0000002e0000002e0000002e0000002e", 7552=>X"0000002e0000002e0000002e0000002e", 7553=>X"0000002e0000002e0000002e0000002e", 7554=>X"0000002e0000002e0000002e0000002e", 
7555=>X"0000002e0000002e0000002e0000002e", 7556=>X"0000002e0000002e0000002e0000002e", 7557=>X"0000002e0000002e0000002e0000002e", 7558=>X"0000002e0000002e0000002e0000002e", 7559=>X"0000002e0000002e0000002e0000002e", 
7560=>X"0000002e0000002e0000002e0000002e", 7561=>X"0000002e0000002e0000002e0000002e", 7562=>X"0000002e0000002e0000002e0000002e", 7563=>X"0000002e0000002e0000002e0000002e", 7564=>X"0000002e0000002e0000002e0000002e", 
7565=>X"0000002e0000002e0000002e0000002e", 7566=>X"0000002e0000002e0000002e0000002e", 7567=>X"0000002e0000002e0000002e0000002e", 7568=>X"0000002e0000002e0000002e0000002e", 7569=>X"0000002e0000002e0000002e0000002e", 
7570=>X"0000002e0000002e0000002e0000002e", 7571=>X"0000002e0000002e0000002e0000002e", 7572=>X"0000002e0000002e0000002e0000002e", 7573=>X"0000002e0000002e0000002e0000002e", 7574=>X"0000002e0000002e0000002e0000002e", 
7575=>X"0000002e0000002e0000002e0000002e", 7576=>X"0000002e0000002e0000002e0000002e", 7577=>X"0000002e0000002e0000002e0000002e", 7578=>X"0000002e0000002e0000002e0000002e", 7579=>X"0000002e0000002e0000002e0000002e", 
7580=>X"0000002e0000002e0000002e0000002e", 7581=>X"0000002e0000002e0000002e0000002e", 7582=>X"0000002e0000002e0000002e0000002e", 7583=>X"0000002e0000002e0000002e0000002e", 7584=>X"0000002e0000002e0000002e0000002e", 
7585=>X"0000002e0000002e0000002e0000002e", 7586=>X"0000002e0000002e0000002e0000002e", 7587=>X"0000002e0000002e0000002e0000002e", 7588=>X"0000002e0000002e0000002e0000002e", 7589=>X"0000002e0000002e0000002e0000002e", 
7590=>X"0000002e0000002e0000002e0000002e", 7591=>X"0000002e0000002e0000002e0000002e", 7592=>X"0000002e0000002e0000002e0000002e", 7593=>X"0000002e0000002e0000002e0000002e", 7594=>X"0000002e0000002e0000002e0000002e", 
7595=>X"0000002e0000002e0000002e0000002e", 7596=>X"0000002e0000002e0000002e0000002e", 7597=>X"0000002e0000002e0000002e0000002e", 7598=>X"0000002e0000002e0000002e0000002e", 7599=>X"0000002e0000002e0000002e0000002e", 
7600=>X"0000002e0000002e0000002e0000002e", 7601=>X"0000002e0000002e0000002e0000002e", 7602=>X"0000002e0000002e0000002e0000002e", 7603=>X"0000002e0000002e0000002e0000002e", 7604=>X"0000002e0000002e0000002e0000002e", 
7605=>X"0000002e0000002e0000002e0000002e", 7606=>X"0000002e0000002e0000002e0000002e", 7607=>X"0000002e0000002e0000002e0000002e", 7608=>X"0000002e0000002e0000002e0000002e", 7609=>X"0000002e0000002e0000002e0000002e", 
7610=>X"0000002e0000002e0000002e0000002e", 7611=>X"0000002e0000002e0000002e0000002e", 7612=>X"0000002e0000002e0000002e0000002e", 7613=>X"0000002e0000002e0000002e0000002e", 7614=>X"0000002e0000002e0000002e0000002e", 
7615=>X"0000002e0000002e0000002e0000002e", 7616=>X"0000002e0000002e0000002e0000002e", 7617=>X"0000002e0000002e0000002e0000002e", 7618=>X"0000002e0000002e0000002e0000002e", 7619=>X"0000002e0000002e0000002e0000002e", 
7620=>X"0000002e0000002e0000002e0000002e", 7621=>X"0000002e0000002e0000002e0000002e", 7622=>X"0000002e0000002e0000002e0000002e", 7623=>X"0000002e0000002e0000002e0000002e", 7624=>X"0000002e0000002e0000002e0000002e", 
7625=>X"0000002e0000002e0000002e0000002e", 7626=>X"0000002e0000002e0000002e0000002e", 7627=>X"0000002e0000002e0000002e0000002e", 7628=>X"0000002e0000002e0000002e0000002e", 7629=>X"0000002e0000002e0000002e0000002e", 
7630=>X"0000002e0000002e0000002e0000002e", 7631=>X"0000002d0000002d0000002d0000002e", 7632=>X"0000002d0000002d0000002d0000002d", 7633=>X"0000002d0000002d0000002d0000002d", 7634=>X"0000002d0000002d0000002d0000002d", 
7635=>X"0000002d0000002d0000002d0000002d", 7636=>X"0000002d0000002d0000002d0000002d", 7637=>X"0000002d0000002d0000002d0000002d", 7638=>X"0000002d0000002d0000002d0000002d", 7639=>X"0000002d0000002d0000002d0000002d", 
7640=>X"0000002d0000002d0000002d0000002d", 7641=>X"0000002d0000002d0000002d0000002d", 7642=>X"0000002d0000002d0000002d0000002d", 7643=>X"0000002d0000002d0000002d0000002d", 7644=>X"0000002d0000002d0000002d0000002d", 
7645=>X"0000002d0000002d0000002d0000002d", 7646=>X"0000002d0000002d0000002d0000002d", 7647=>X"0000002d0000002d0000002d0000002d", 7648=>X"0000002d0000002d0000002d0000002d", 7649=>X"0000002d0000002d0000002d0000002d", 
7650=>X"0000002d0000002d0000002d0000002d", 7651=>X"0000002d0000002d0000002d0000002d", 7652=>X"0000002d0000002d0000002d0000002d", 7653=>X"0000002d0000002d0000002d0000002d", 7654=>X"0000002d0000002d0000002d0000002d", 
7655=>X"0000002d0000002d0000002d0000002d", 7656=>X"0000002d0000002d0000002d0000002d", 7657=>X"0000002d0000002d0000002d0000002d", 7658=>X"0000002d0000002d0000002d0000002d", 7659=>X"0000002d0000002d0000002d0000002d", 
7660=>X"0000002d0000002d0000002d0000002d", 7661=>X"0000002d0000002d0000002d0000002d", 7662=>X"0000002d0000002d0000002d0000002d", 7663=>X"0000002d0000002d0000002d0000002d", 7664=>X"0000002d0000002d0000002d0000002d", 
7665=>X"0000002d0000002d0000002d0000002d", 7666=>X"0000002d0000002d0000002d0000002d", 7667=>X"0000002d0000002d0000002d0000002d", 7668=>X"0000002d0000002d0000002d0000002d", 7669=>X"0000002d0000002d0000002d0000002d", 
7670=>X"0000002d0000002d0000002d0000002d", 7671=>X"0000002d0000002d0000002d0000002d", 7672=>X"0000002d0000002d0000002d0000002d", 7673=>X"0000002d0000002d0000002d0000002d", 7674=>X"0000002d0000002d0000002d0000002d", 
7675=>X"0000002d0000002d0000002d0000002d", 7676=>X"0000002d0000002d0000002d0000002d", 7677=>X"0000002d0000002d0000002d0000002d", 7678=>X"0000002d0000002d0000002d0000002d", 7679=>X"0000002d0000002d0000002d0000002d", 
7680=>X"0000002d0000002d0000002d0000002d", 7681=>X"0000002d0000002d0000002d0000002d", 7682=>X"0000002d0000002d0000002d0000002d", 7683=>X"0000002d0000002d0000002d0000002d", 7684=>X"0000002d0000002d0000002d0000002d", 
7685=>X"0000002d0000002d0000002d0000002d", 7686=>X"0000002d0000002d0000002d0000002d", 7687=>X"0000002d0000002d0000002d0000002d", 7688=>X"0000002d0000002d0000002d0000002d", 7689=>X"0000002d0000002d0000002d0000002d", 
7690=>X"0000002d0000002d0000002d0000002d", 7691=>X"0000002d0000002d0000002d0000002d", 7692=>X"0000002d0000002d0000002d0000002d", 7693=>X"0000002d0000002d0000002d0000002d", 7694=>X"0000002d0000002d0000002d0000002d", 
7695=>X"0000002d0000002d0000002d0000002d", 7696=>X"0000002d0000002d0000002d0000002d", 7697=>X"0000002d0000002d0000002d0000002d", 7698=>X"0000002d0000002d0000002d0000002d", 7699=>X"0000002d0000002d0000002d0000002d", 
7700=>X"0000002d0000002d0000002d0000002d", 7701=>X"0000002d0000002d0000002d0000002d", 7702=>X"0000002d0000002d0000002d0000002d", 7703=>X"0000002d0000002d0000002d0000002d", 7704=>X"0000002d0000002d0000002d0000002d", 
7705=>X"0000002d0000002d0000002d0000002d", 7706=>X"0000002d0000002d0000002d0000002d", 7707=>X"0000002d0000002d0000002d0000002d", 7708=>X"0000002d0000002d0000002d0000002d", 7709=>X"0000002d0000002d0000002d0000002d", 
7710=>X"0000002d0000002d0000002d0000002d", 7711=>X"0000002d0000002d0000002d0000002d", 7712=>X"0000002d0000002d0000002d0000002d", 7713=>X"0000002d0000002d0000002d0000002d", 7714=>X"0000002d0000002d0000002d0000002d", 
7715=>X"0000002d0000002d0000002d0000002d", 7716=>X"0000002d0000002d0000002d0000002d", 7717=>X"0000002d0000002d0000002d0000002d", 7718=>X"0000002d0000002d0000002d0000002d", 7719=>X"0000002d0000002d0000002d0000002d", 
7720=>X"0000002d0000002d0000002d0000002d", 7721=>X"0000002d0000002d0000002d0000002d", 7722=>X"0000002d0000002d0000002d0000002d", 7723=>X"0000002d0000002d0000002d0000002d", 7724=>X"0000002d0000002d0000002d0000002d", 
7725=>X"0000002d0000002d0000002d0000002d", 7726=>X"0000002d0000002d0000002d0000002d", 7727=>X"0000002d0000002d0000002d0000002d", 7728=>X"0000002d0000002d0000002d0000002d", 7729=>X"0000002d0000002d0000002d0000002d", 
7730=>X"0000002d0000002d0000002d0000002d", 7731=>X"0000002d0000002d0000002d0000002d", 7732=>X"0000002d0000002d0000002d0000002d", 7733=>X"0000002d0000002d0000002d0000002d", 7734=>X"0000002d0000002d0000002d0000002d", 
7735=>X"0000002d0000002d0000002d0000002d", 7736=>X"0000002d0000002d0000002d0000002d", 7737=>X"0000002d0000002d0000002d0000002d", 7738=>X"0000002d0000002d0000002d0000002d", 7739=>X"0000002d0000002d0000002d0000002d", 
7740=>X"0000002d0000002d0000002d0000002d", 7741=>X"0000002d0000002d0000002d0000002d", 7742=>X"0000002d0000002d0000002d0000002d", 7743=>X"0000002d0000002d0000002d0000002d", 7744=>X"0000002d0000002d0000002d0000002d", 
7745=>X"0000002d0000002d0000002d0000002d", 7746=>X"0000002d0000002d0000002d0000002d", 7747=>X"0000002d0000002d0000002d0000002d", 7748=>X"0000002d0000002d0000002d0000002d", 7749=>X"0000002d0000002d0000002d0000002d", 
7750=>X"0000002d0000002d0000002d0000002d", 7751=>X"0000002d0000002d0000002d0000002d", 7752=>X"0000002d0000002d0000002d0000002d", 7753=>X"0000002d0000002d0000002d0000002d", 7754=>X"0000002d0000002d0000002d0000002d", 
7755=>X"0000002d0000002d0000002d0000002d", 7756=>X"0000002d0000002d0000002d0000002d", 7757=>X"0000002d0000002d0000002d0000002d", 7758=>X"0000002d0000002d0000002d0000002d", 7759=>X"0000002d0000002d0000002d0000002d", 
7760=>X"0000002c0000002d0000002d0000002d", 7761=>X"0000002c0000002c0000002c0000002c", 7762=>X"0000002c0000002c0000002c0000002c", 7763=>X"0000002c0000002c0000002c0000002c", 7764=>X"0000002c0000002c0000002c0000002c", 
7765=>X"0000002c0000002c0000002c0000002c", 7766=>X"0000002c0000002c0000002c0000002c", 7767=>X"0000002c0000002c0000002c0000002c", 7768=>X"0000002c0000002c0000002c0000002c", 7769=>X"0000002c0000002c0000002c0000002c", 
7770=>X"0000002c0000002c0000002c0000002c", 7771=>X"0000002c0000002c0000002c0000002c", 7772=>X"0000002c0000002c0000002c0000002c", 7773=>X"0000002c0000002c0000002c0000002c", 7774=>X"0000002c0000002c0000002c0000002c", 
7775=>X"0000002c0000002c0000002c0000002c", 7776=>X"0000002c0000002c0000002c0000002c", 7777=>X"0000002c0000002c0000002c0000002c", 7778=>X"0000002c0000002c0000002c0000002c", 7779=>X"0000002c0000002c0000002c0000002c", 
7780=>X"0000002c0000002c0000002c0000002c", 7781=>X"0000002c0000002c0000002c0000002c", 7782=>X"0000002c0000002c0000002c0000002c", 7783=>X"0000002c0000002c0000002c0000002c", 7784=>X"0000002c0000002c0000002c0000002c", 
7785=>X"0000002c0000002c0000002c0000002c", 7786=>X"0000002c0000002c0000002c0000002c", 7787=>X"0000002c0000002c0000002c0000002c", 7788=>X"0000002c0000002c0000002c0000002c", 7789=>X"0000002c0000002c0000002c0000002c", 
7790=>X"0000002c0000002c0000002c0000002c", 7791=>X"0000002c0000002c0000002c0000002c", 7792=>X"0000002c0000002c0000002c0000002c", 7793=>X"0000002c0000002c0000002c0000002c", 7794=>X"0000002c0000002c0000002c0000002c", 
7795=>X"0000002c0000002c0000002c0000002c", 7796=>X"0000002c0000002c0000002c0000002c", 7797=>X"0000002c0000002c0000002c0000002c", 7798=>X"0000002c0000002c0000002c0000002c", 7799=>X"0000002c0000002c0000002c0000002c", 
7800=>X"0000002c0000002c0000002c0000002c", 7801=>X"0000002c0000002c0000002c0000002c", 7802=>X"0000002c0000002c0000002c0000002c", 7803=>X"0000002c0000002c0000002c0000002c", 7804=>X"0000002c0000002c0000002c0000002c", 
7805=>X"0000002c0000002c0000002c0000002c", 7806=>X"0000002c0000002c0000002c0000002c", 7807=>X"0000002c0000002c0000002c0000002c", 7808=>X"0000002c0000002c0000002c0000002c", 7809=>X"0000002c0000002c0000002c0000002c", 
7810=>X"0000002c0000002c0000002c0000002c", 7811=>X"0000002c0000002c0000002c0000002c", 7812=>X"0000002c0000002c0000002c0000002c", 7813=>X"0000002c0000002c0000002c0000002c", 7814=>X"0000002c0000002c0000002c0000002c", 
7815=>X"0000002c0000002c0000002c0000002c", 7816=>X"0000002c0000002c0000002c0000002c", 7817=>X"0000002c0000002c0000002c0000002c", 7818=>X"0000002c0000002c0000002c0000002c", 7819=>X"0000002c0000002c0000002c0000002c", 
7820=>X"0000002c0000002c0000002c0000002c", 7821=>X"0000002c0000002c0000002c0000002c", 7822=>X"0000002c0000002c0000002c0000002c", 7823=>X"0000002c0000002c0000002c0000002c", 7824=>X"0000002c0000002c0000002c0000002c", 
7825=>X"0000002c0000002c0000002c0000002c", 7826=>X"0000002c0000002c0000002c0000002c", 7827=>X"0000002c0000002c0000002c0000002c", 7828=>X"0000002c0000002c0000002c0000002c", 7829=>X"0000002c0000002c0000002c0000002c", 
7830=>X"0000002c0000002c0000002c0000002c", 7831=>X"0000002c0000002c0000002c0000002c", 7832=>X"0000002c0000002c0000002c0000002c", 7833=>X"0000002c0000002c0000002c0000002c", 7834=>X"0000002c0000002c0000002c0000002c", 
7835=>X"0000002c0000002c0000002c0000002c", 7836=>X"0000002c0000002c0000002c0000002c", 7837=>X"0000002c0000002c0000002c0000002c", 7838=>X"0000002c0000002c0000002c0000002c", 7839=>X"0000002c0000002c0000002c0000002c", 
7840=>X"0000002c0000002c0000002c0000002c", 7841=>X"0000002c0000002c0000002c0000002c", 7842=>X"0000002c0000002c0000002c0000002c", 7843=>X"0000002c0000002c0000002c0000002c", 7844=>X"0000002c0000002c0000002c0000002c", 
7845=>X"0000002c0000002c0000002c0000002c", 7846=>X"0000002c0000002c0000002c0000002c", 7847=>X"0000002c0000002c0000002c0000002c", 7848=>X"0000002c0000002c0000002c0000002c", 7849=>X"0000002c0000002c0000002c0000002c", 
7850=>X"0000002c0000002c0000002c0000002c", 7851=>X"0000002c0000002c0000002c0000002c", 7852=>X"0000002c0000002c0000002c0000002c", 7853=>X"0000002c0000002c0000002c0000002c", 7854=>X"0000002c0000002c0000002c0000002c", 
7855=>X"0000002c0000002c0000002c0000002c", 7856=>X"0000002c0000002c0000002c0000002c", 7857=>X"0000002c0000002c0000002c0000002c", 7858=>X"0000002c0000002c0000002c0000002c", 7859=>X"0000002c0000002c0000002c0000002c", 
7860=>X"0000002c0000002c0000002c0000002c", 7861=>X"0000002c0000002c0000002c0000002c", 7862=>X"0000002c0000002c0000002c0000002c", 7863=>X"0000002c0000002c0000002c0000002c", 7864=>X"0000002c0000002c0000002c0000002c", 
7865=>X"0000002c0000002c0000002c0000002c", 7866=>X"0000002c0000002c0000002c0000002c", 7867=>X"0000002c0000002c0000002c0000002c", 7868=>X"0000002c0000002c0000002c0000002c", 7869=>X"0000002c0000002c0000002c0000002c", 
7870=>X"0000002c0000002c0000002c0000002c", 7871=>X"0000002c0000002c0000002c0000002c", 7872=>X"0000002c0000002c0000002c0000002c", 7873=>X"0000002c0000002c0000002c0000002c", 7874=>X"0000002c0000002c0000002c0000002c", 
7875=>X"0000002c0000002c0000002c0000002c", 7876=>X"0000002c0000002c0000002c0000002c", 7877=>X"0000002c0000002c0000002c0000002c", 7878=>X"0000002c0000002c0000002c0000002c", 7879=>X"0000002c0000002c0000002c0000002c", 
7880=>X"0000002c0000002c0000002c0000002c", 7881=>X"0000002c0000002c0000002c0000002c", 7882=>X"0000002c0000002c0000002c0000002c", 7883=>X"0000002c0000002c0000002c0000002c", 7884=>X"0000002c0000002c0000002c0000002c", 
7885=>X"0000002c0000002c0000002c0000002c", 7886=>X"0000002c0000002c0000002c0000002c", 7887=>X"0000002c0000002c0000002c0000002c", 7888=>X"0000002c0000002c0000002c0000002c", 7889=>X"0000002c0000002c0000002c0000002c", 
7890=>X"0000002c0000002c0000002c0000002c", 7891=>X"0000002c0000002c0000002c0000002c", 7892=>X"0000002c0000002c0000002c0000002c", 7893=>X"0000002c0000002c0000002c0000002c", 7894=>X"0000002c0000002c0000002c0000002c", 
7895=>X"0000002c0000002c0000002c0000002c", 7896=>X"0000002b0000002b0000002b0000002c", 7897=>X"0000002b0000002b0000002b0000002b", 7898=>X"0000002b0000002b0000002b0000002b", 7899=>X"0000002b0000002b0000002b0000002b", 
7900=>X"0000002b0000002b0000002b0000002b", 7901=>X"0000002b0000002b0000002b0000002b", 7902=>X"0000002b0000002b0000002b0000002b", 7903=>X"0000002b0000002b0000002b0000002b", 7904=>X"0000002b0000002b0000002b0000002b", 
7905=>X"0000002b0000002b0000002b0000002b", 7906=>X"0000002b0000002b0000002b0000002b", 7907=>X"0000002b0000002b0000002b0000002b", 7908=>X"0000002b0000002b0000002b0000002b", 7909=>X"0000002b0000002b0000002b0000002b", 
7910=>X"0000002b0000002b0000002b0000002b", 7911=>X"0000002b0000002b0000002b0000002b", 7912=>X"0000002b0000002b0000002b0000002b", 7913=>X"0000002b0000002b0000002b0000002b", 7914=>X"0000002b0000002b0000002b0000002b", 
7915=>X"0000002b0000002b0000002b0000002b", 7916=>X"0000002b0000002b0000002b0000002b", 7917=>X"0000002b0000002b0000002b0000002b", 7918=>X"0000002b0000002b0000002b0000002b", 7919=>X"0000002b0000002b0000002b0000002b", 
7920=>X"0000002b0000002b0000002b0000002b", 7921=>X"0000002b0000002b0000002b0000002b", 7922=>X"0000002b0000002b0000002b0000002b", 7923=>X"0000002b0000002b0000002b0000002b", 7924=>X"0000002b0000002b0000002b0000002b", 
7925=>X"0000002b0000002b0000002b0000002b", 7926=>X"0000002b0000002b0000002b0000002b", 7927=>X"0000002b0000002b0000002b0000002b", 7928=>X"0000002b0000002b0000002b0000002b", 7929=>X"0000002b0000002b0000002b0000002b", 
7930=>X"0000002b0000002b0000002b0000002b", 7931=>X"0000002b0000002b0000002b0000002b", 7932=>X"0000002b0000002b0000002b0000002b", 7933=>X"0000002b0000002b0000002b0000002b", 7934=>X"0000002b0000002b0000002b0000002b", 
7935=>X"0000002b0000002b0000002b0000002b", 7936=>X"0000002b0000002b0000002b0000002b", 7937=>X"0000002b0000002b0000002b0000002b", 7938=>X"0000002b0000002b0000002b0000002b", 7939=>X"0000002b0000002b0000002b0000002b", 
7940=>X"0000002b0000002b0000002b0000002b", 7941=>X"0000002b0000002b0000002b0000002b", 7942=>X"0000002b0000002b0000002b0000002b", 7943=>X"0000002b0000002b0000002b0000002b", 7944=>X"0000002b0000002b0000002b0000002b", 
7945=>X"0000002b0000002b0000002b0000002b", 7946=>X"0000002b0000002b0000002b0000002b", 7947=>X"0000002b0000002b0000002b0000002b", 7948=>X"0000002b0000002b0000002b0000002b", 7949=>X"0000002b0000002b0000002b0000002b", 
7950=>X"0000002b0000002b0000002b0000002b", 7951=>X"0000002b0000002b0000002b0000002b", 7952=>X"0000002b0000002b0000002b0000002b", 7953=>X"0000002b0000002b0000002b0000002b", 7954=>X"0000002b0000002b0000002b0000002b", 
7955=>X"0000002b0000002b0000002b0000002b", 7956=>X"0000002b0000002b0000002b0000002b", 7957=>X"0000002b0000002b0000002b0000002b", 7958=>X"0000002b0000002b0000002b0000002b", 7959=>X"0000002b0000002b0000002b0000002b", 
7960=>X"0000002b0000002b0000002b0000002b", 7961=>X"0000002b0000002b0000002b0000002b", 7962=>X"0000002b0000002b0000002b0000002b", 7963=>X"0000002b0000002b0000002b0000002b", 7964=>X"0000002b0000002b0000002b0000002b", 
7965=>X"0000002b0000002b0000002b0000002b", 7966=>X"0000002b0000002b0000002b0000002b", 7967=>X"0000002b0000002b0000002b0000002b", 7968=>X"0000002b0000002b0000002b0000002b", 7969=>X"0000002b0000002b0000002b0000002b", 
7970=>X"0000002b0000002b0000002b0000002b", 7971=>X"0000002b0000002b0000002b0000002b", 7972=>X"0000002b0000002b0000002b0000002b", 7973=>X"0000002b0000002b0000002b0000002b", 7974=>X"0000002b0000002b0000002b0000002b", 
7975=>X"0000002b0000002b0000002b0000002b", 7976=>X"0000002b0000002b0000002b0000002b", 7977=>X"0000002b0000002b0000002b0000002b", 7978=>X"0000002b0000002b0000002b0000002b", 7979=>X"0000002b0000002b0000002b0000002b", 
7980=>X"0000002b0000002b0000002b0000002b", 7981=>X"0000002b0000002b0000002b0000002b", 7982=>X"0000002b0000002b0000002b0000002b", 7983=>X"0000002b0000002b0000002b0000002b", 7984=>X"0000002b0000002b0000002b0000002b", 
7985=>X"0000002b0000002b0000002b0000002b", 7986=>X"0000002b0000002b0000002b0000002b", 7987=>X"0000002b0000002b0000002b0000002b", 7988=>X"0000002b0000002b0000002b0000002b", 7989=>X"0000002b0000002b0000002b0000002b", 
7990=>X"0000002b0000002b0000002b0000002b", 7991=>X"0000002b0000002b0000002b0000002b", 7992=>X"0000002b0000002b0000002b0000002b", 7993=>X"0000002b0000002b0000002b0000002b", 7994=>X"0000002b0000002b0000002b0000002b", 
7995=>X"0000002b0000002b0000002b0000002b", 7996=>X"0000002b0000002b0000002b0000002b", 7997=>X"0000002b0000002b0000002b0000002b", 7998=>X"0000002b0000002b0000002b0000002b", 7999=>X"0000002b0000002b0000002b0000002b", 
8000=>X"0000002b0000002b0000002b0000002b", 8001=>X"0000002b0000002b0000002b0000002b", 8002=>X"0000002b0000002b0000002b0000002b", 8003=>X"0000002b0000002b0000002b0000002b", 8004=>X"0000002b0000002b0000002b0000002b", 
8005=>X"0000002b0000002b0000002b0000002b", 8006=>X"0000002b0000002b0000002b0000002b", 8007=>X"0000002b0000002b0000002b0000002b", 8008=>X"0000002b0000002b0000002b0000002b", 8009=>X"0000002b0000002b0000002b0000002b", 
8010=>X"0000002b0000002b0000002b0000002b", 8011=>X"0000002b0000002b0000002b0000002b", 8012=>X"0000002b0000002b0000002b0000002b", 8013=>X"0000002b0000002b0000002b0000002b", 8014=>X"0000002b0000002b0000002b0000002b", 
8015=>X"0000002b0000002b0000002b0000002b", 8016=>X"0000002b0000002b0000002b0000002b", 8017=>X"0000002b0000002b0000002b0000002b", 8018=>X"0000002b0000002b0000002b0000002b", 8019=>X"0000002b0000002b0000002b0000002b", 
8020=>X"0000002b0000002b0000002b0000002b", 8021=>X"0000002b0000002b0000002b0000002b", 8022=>X"0000002b0000002b0000002b0000002b", 8023=>X"0000002b0000002b0000002b0000002b", 8024=>X"0000002b0000002b0000002b0000002b", 
8025=>X"0000002b0000002b0000002b0000002b", 8026=>X"0000002b0000002b0000002b0000002b", 8027=>X"0000002b0000002b0000002b0000002b", 8028=>X"0000002b0000002b0000002b0000002b", 8029=>X"0000002b0000002b0000002b0000002b", 
8030=>X"0000002b0000002b0000002b0000002b", 8031=>X"0000002b0000002b0000002b0000002b", 8032=>X"0000002b0000002b0000002b0000002b", 8033=>X"0000002b0000002b0000002b0000002b", 8034=>X"0000002b0000002b0000002b0000002b", 
8035=>X"0000002b0000002b0000002b0000002b", 8036=>X"0000002b0000002b0000002b0000002b", 8037=>X"0000002b0000002b0000002b0000002b", 8038=>X"0000002a0000002a0000002a0000002a", 8039=>X"0000002a0000002a0000002a0000002a", 
8040=>X"0000002a0000002a0000002a0000002a", 8041=>X"0000002a0000002a0000002a0000002a", 8042=>X"0000002a0000002a0000002a0000002a", 8043=>X"0000002a0000002a0000002a0000002a", 8044=>X"0000002a0000002a0000002a0000002a", 
8045=>X"0000002a0000002a0000002a0000002a", 8046=>X"0000002a0000002a0000002a0000002a", 8047=>X"0000002a0000002a0000002a0000002a", 8048=>X"0000002a0000002a0000002a0000002a", 8049=>X"0000002a0000002a0000002a0000002a", 
8050=>X"0000002a0000002a0000002a0000002a", 8051=>X"0000002a0000002a0000002a0000002a", 8052=>X"0000002a0000002a0000002a0000002a", 8053=>X"0000002a0000002a0000002a0000002a", 8054=>X"0000002a0000002a0000002a0000002a", 
8055=>X"0000002a0000002a0000002a0000002a", 8056=>X"0000002a0000002a0000002a0000002a", 8057=>X"0000002a0000002a0000002a0000002a", 8058=>X"0000002a0000002a0000002a0000002a", 8059=>X"0000002a0000002a0000002a0000002a", 
8060=>X"0000002a0000002a0000002a0000002a", 8061=>X"0000002a0000002a0000002a0000002a", 8062=>X"0000002a0000002a0000002a0000002a", 8063=>X"0000002a0000002a0000002a0000002a", 8064=>X"0000002a0000002a0000002a0000002a", 
8065=>X"0000002a0000002a0000002a0000002a", 8066=>X"0000002a0000002a0000002a0000002a", 8067=>X"0000002a0000002a0000002a0000002a", 8068=>X"0000002a0000002a0000002a0000002a", 8069=>X"0000002a0000002a0000002a0000002a", 
8070=>X"0000002a0000002a0000002a0000002a", 8071=>X"0000002a0000002a0000002a0000002a", 8072=>X"0000002a0000002a0000002a0000002a", 8073=>X"0000002a0000002a0000002a0000002a", 8074=>X"0000002a0000002a0000002a0000002a", 
8075=>X"0000002a0000002a0000002a0000002a", 8076=>X"0000002a0000002a0000002a0000002a", 8077=>X"0000002a0000002a0000002a0000002a", 8078=>X"0000002a0000002a0000002a0000002a", 8079=>X"0000002a0000002a0000002a0000002a", 
8080=>X"0000002a0000002a0000002a0000002a", 8081=>X"0000002a0000002a0000002a0000002a", 8082=>X"0000002a0000002a0000002a0000002a", 8083=>X"0000002a0000002a0000002a0000002a", 8084=>X"0000002a0000002a0000002a0000002a", 
8085=>X"0000002a0000002a0000002a0000002a", 8086=>X"0000002a0000002a0000002a0000002a", 8087=>X"0000002a0000002a0000002a0000002a", 8088=>X"0000002a0000002a0000002a0000002a", 8089=>X"0000002a0000002a0000002a0000002a", 
8090=>X"0000002a0000002a0000002a0000002a", 8091=>X"0000002a0000002a0000002a0000002a", 8092=>X"0000002a0000002a0000002a0000002a", 8093=>X"0000002a0000002a0000002a0000002a", 8094=>X"0000002a0000002a0000002a0000002a", 
8095=>X"0000002a0000002a0000002a0000002a", 8096=>X"0000002a0000002a0000002a0000002a", 8097=>X"0000002a0000002a0000002a0000002a", 8098=>X"0000002a0000002a0000002a0000002a", 8099=>X"0000002a0000002a0000002a0000002a", 
8100=>X"0000002a0000002a0000002a0000002a", 8101=>X"0000002a0000002a0000002a0000002a", 8102=>X"0000002a0000002a0000002a0000002a", 8103=>X"0000002a0000002a0000002a0000002a", 8104=>X"0000002a0000002a0000002a0000002a", 
8105=>X"0000002a0000002a0000002a0000002a", 8106=>X"0000002a0000002a0000002a0000002a", 8107=>X"0000002a0000002a0000002a0000002a", 8108=>X"0000002a0000002a0000002a0000002a", 8109=>X"0000002a0000002a0000002a0000002a", 
8110=>X"0000002a0000002a0000002a0000002a", 8111=>X"0000002a0000002a0000002a0000002a", 8112=>X"0000002a0000002a0000002a0000002a", 8113=>X"0000002a0000002a0000002a0000002a", 8114=>X"0000002a0000002a0000002a0000002a", 
8115=>X"0000002a0000002a0000002a0000002a", 8116=>X"0000002a0000002a0000002a0000002a", 8117=>X"0000002a0000002a0000002a0000002a", 8118=>X"0000002a0000002a0000002a0000002a", 8119=>X"0000002a0000002a0000002a0000002a", 
8120=>X"0000002a0000002a0000002a0000002a", 8121=>X"0000002a0000002a0000002a0000002a", 8122=>X"0000002a0000002a0000002a0000002a", 8123=>X"0000002a0000002a0000002a0000002a", 8124=>X"0000002a0000002a0000002a0000002a", 
8125=>X"0000002a0000002a0000002a0000002a", 8126=>X"0000002a0000002a0000002a0000002a", 8127=>X"0000002a0000002a0000002a0000002a", 8128=>X"0000002a0000002a0000002a0000002a", 8129=>X"0000002a0000002a0000002a0000002a", 
8130=>X"0000002a0000002a0000002a0000002a", 8131=>X"0000002a0000002a0000002a0000002a", 8132=>X"0000002a0000002a0000002a0000002a", 8133=>X"0000002a0000002a0000002a0000002a", 8134=>X"0000002a0000002a0000002a0000002a", 
8135=>X"0000002a0000002a0000002a0000002a", 8136=>X"0000002a0000002a0000002a0000002a", 8137=>X"0000002a0000002a0000002a0000002a", 8138=>X"0000002a0000002a0000002a0000002a", 8139=>X"0000002a0000002a0000002a0000002a", 
8140=>X"0000002a0000002a0000002a0000002a", 8141=>X"0000002a0000002a0000002a0000002a", 8142=>X"0000002a0000002a0000002a0000002a", 8143=>X"0000002a0000002a0000002a0000002a", 8144=>X"0000002a0000002a0000002a0000002a", 
8145=>X"0000002a0000002a0000002a0000002a", 8146=>X"0000002a0000002a0000002a0000002a", 8147=>X"0000002a0000002a0000002a0000002a", 8148=>X"0000002a0000002a0000002a0000002a", 8149=>X"0000002a0000002a0000002a0000002a", 
8150=>X"0000002a0000002a0000002a0000002a", 8151=>X"0000002a0000002a0000002a0000002a", 8152=>X"0000002a0000002a0000002a0000002a", 8153=>X"0000002a0000002a0000002a0000002a", 8154=>X"0000002a0000002a0000002a0000002a", 
8155=>X"0000002a0000002a0000002a0000002a", 8156=>X"0000002a0000002a0000002a0000002a", 8157=>X"0000002a0000002a0000002a0000002a", 8158=>X"0000002a0000002a0000002a0000002a", 8159=>X"0000002a0000002a0000002a0000002a", 
8160=>X"0000002a0000002a0000002a0000002a", 8161=>X"0000002a0000002a0000002a0000002a", 8162=>X"0000002a0000002a0000002a0000002a", 8163=>X"0000002a0000002a0000002a0000002a", 8164=>X"0000002a0000002a0000002a0000002a", 
8165=>X"0000002a0000002a0000002a0000002a", 8166=>X"0000002a0000002a0000002a0000002a", 8167=>X"0000002a0000002a0000002a0000002a", 8168=>X"0000002a0000002a0000002a0000002a", 8169=>X"0000002a0000002a0000002a0000002a", 
8170=>X"0000002a0000002a0000002a0000002a", 8171=>X"0000002a0000002a0000002a0000002a", 8172=>X"0000002a0000002a0000002a0000002a", 8173=>X"0000002a0000002a0000002a0000002a", 8174=>X"0000002a0000002a0000002a0000002a", 
8175=>X"0000002a0000002a0000002a0000002a", 8176=>X"0000002a0000002a0000002a0000002a", 8177=>X"0000002a0000002a0000002a0000002a", 8178=>X"0000002a0000002a0000002a0000002a", 8179=>X"0000002a0000002a0000002a0000002a", 
8180=>X"0000002a0000002a0000002a0000002a", 8181=>X"0000002a0000002a0000002a0000002a", 8182=>X"0000002a0000002a0000002a0000002a", 8183=>X"0000002a0000002a0000002a0000002a", 8184=>X"0000002a0000002a0000002a0000002a", 
8185=>X"0000002a0000002a0000002a0000002a", 8186=>X"00000029000000290000002a0000002a", 8187=>X"00000029000000290000002900000029", 8188=>X"00000029000000290000002900000029", 8189=>X"00000029000000290000002900000029", 
8190=>X"00000029000000290000002900000029", 8191=>X"00000029000000290000002900000029", 8192=>X"00000029000000290000002900000029", 8193=>X"00000029000000290000002900000029", 8194=>X"00000029000000290000002900000029", 
8195=>X"00000029000000290000002900000029", 8196=>X"00000029000000290000002900000029", 8197=>X"00000029000000290000002900000029", 8198=>X"00000029000000290000002900000029", 8199=>X"00000029000000290000002900000029", 
8200=>X"00000029000000290000002900000029", 8201=>X"00000029000000290000002900000029", 8202=>X"00000029000000290000002900000029", 8203=>X"00000029000000290000002900000029", 8204=>X"00000029000000290000002900000029", 
8205=>X"00000029000000290000002900000029", 8206=>X"00000029000000290000002900000029", 8207=>X"00000029000000290000002900000029", 8208=>X"00000029000000290000002900000029", 8209=>X"00000029000000290000002900000029", 
8210=>X"00000029000000290000002900000029", 8211=>X"00000029000000290000002900000029", 8212=>X"00000029000000290000002900000029", 8213=>X"00000029000000290000002900000029", 8214=>X"00000029000000290000002900000029", 
8215=>X"00000029000000290000002900000029", 8216=>X"00000029000000290000002900000029", 8217=>X"00000029000000290000002900000029", 8218=>X"00000029000000290000002900000029", 8219=>X"00000029000000290000002900000029", 
8220=>X"00000029000000290000002900000029", 8221=>X"00000029000000290000002900000029", 8222=>X"00000029000000290000002900000029", 8223=>X"00000029000000290000002900000029", 8224=>X"00000029000000290000002900000029", 
8225=>X"00000029000000290000002900000029", 8226=>X"00000029000000290000002900000029", 8227=>X"00000029000000290000002900000029", 8228=>X"00000029000000290000002900000029", 8229=>X"00000029000000290000002900000029", 
8230=>X"00000029000000290000002900000029", 8231=>X"00000029000000290000002900000029", 8232=>X"00000029000000290000002900000029", 8233=>X"00000029000000290000002900000029", 8234=>X"00000029000000290000002900000029", 
8235=>X"00000029000000290000002900000029", 8236=>X"00000029000000290000002900000029", 8237=>X"00000029000000290000002900000029", 8238=>X"00000029000000290000002900000029", 8239=>X"00000029000000290000002900000029", 
8240=>X"00000029000000290000002900000029", 8241=>X"00000029000000290000002900000029", 8242=>X"00000029000000290000002900000029", 8243=>X"00000029000000290000002900000029", 8244=>X"00000029000000290000002900000029", 
8245=>X"00000029000000290000002900000029", 8246=>X"00000029000000290000002900000029", 8247=>X"00000029000000290000002900000029", 8248=>X"00000029000000290000002900000029", 8249=>X"00000029000000290000002900000029", 
8250=>X"00000029000000290000002900000029", 8251=>X"00000029000000290000002900000029", 8252=>X"00000029000000290000002900000029", 8253=>X"00000029000000290000002900000029", 8254=>X"00000029000000290000002900000029", 
8255=>X"00000029000000290000002900000029", 8256=>X"00000029000000290000002900000029", 8257=>X"00000029000000290000002900000029", 8258=>X"00000029000000290000002900000029", 8259=>X"00000029000000290000002900000029", 
8260=>X"00000029000000290000002900000029", 8261=>X"00000029000000290000002900000029", 8262=>X"00000029000000290000002900000029", 8263=>X"00000029000000290000002900000029", 8264=>X"00000029000000290000002900000029", 
8265=>X"00000029000000290000002900000029", 8266=>X"00000029000000290000002900000029", 8267=>X"00000029000000290000002900000029", 8268=>X"00000029000000290000002900000029", 8269=>X"00000029000000290000002900000029", 
8270=>X"00000029000000290000002900000029", 8271=>X"00000029000000290000002900000029", 8272=>X"00000029000000290000002900000029", 8273=>X"00000029000000290000002900000029", 8274=>X"00000029000000290000002900000029", 
8275=>X"00000029000000290000002900000029", 8276=>X"00000029000000290000002900000029", 8277=>X"00000029000000290000002900000029", 8278=>X"00000029000000290000002900000029", 8279=>X"00000029000000290000002900000029", 
8280=>X"00000029000000290000002900000029", 8281=>X"00000029000000290000002900000029", 8282=>X"00000029000000290000002900000029", 8283=>X"00000029000000290000002900000029", 8284=>X"00000029000000290000002900000029", 
8285=>X"00000029000000290000002900000029", 8286=>X"00000029000000290000002900000029", 8287=>X"00000029000000290000002900000029", 8288=>X"00000029000000290000002900000029", 8289=>X"00000029000000290000002900000029", 
8290=>X"00000029000000290000002900000029", 8291=>X"00000029000000290000002900000029", 8292=>X"00000029000000290000002900000029", 8293=>X"00000029000000290000002900000029", 8294=>X"00000029000000290000002900000029", 
8295=>X"00000029000000290000002900000029", 8296=>X"00000029000000290000002900000029", 8297=>X"00000029000000290000002900000029", 8298=>X"00000029000000290000002900000029", 8299=>X"00000029000000290000002900000029", 
8300=>X"00000029000000290000002900000029", 8301=>X"00000029000000290000002900000029", 8302=>X"00000029000000290000002900000029", 8303=>X"00000029000000290000002900000029", 8304=>X"00000029000000290000002900000029", 
8305=>X"00000029000000290000002900000029", 8306=>X"00000029000000290000002900000029", 8307=>X"00000029000000290000002900000029", 8308=>X"00000029000000290000002900000029", 8309=>X"00000029000000290000002900000029", 
8310=>X"00000029000000290000002900000029", 8311=>X"00000029000000290000002900000029", 8312=>X"00000029000000290000002900000029", 8313=>X"00000029000000290000002900000029", 8314=>X"00000029000000290000002900000029", 
8315=>X"00000029000000290000002900000029", 8316=>X"00000029000000290000002900000029", 8317=>X"00000029000000290000002900000029", 8318=>X"00000029000000290000002900000029", 8319=>X"00000029000000290000002900000029", 
8320=>X"00000029000000290000002900000029", 8321=>X"00000029000000290000002900000029", 8322=>X"00000029000000290000002900000029", 8323=>X"00000029000000290000002900000029", 8324=>X"00000029000000290000002900000029", 
8325=>X"00000029000000290000002900000029", 8326=>X"00000029000000290000002900000029", 8327=>X"00000029000000290000002900000029", 8328=>X"00000029000000290000002900000029", 8329=>X"00000029000000290000002900000029", 
8330=>X"00000029000000290000002900000029", 8331=>X"00000029000000290000002900000029", 8332=>X"00000029000000290000002900000029", 8333=>X"00000029000000290000002900000029", 8334=>X"00000029000000290000002900000029", 
8335=>X"00000029000000290000002900000029", 8336=>X"00000029000000290000002900000029", 8337=>X"00000029000000290000002900000029", 8338=>X"00000029000000290000002900000029", 8339=>X"00000029000000290000002900000029", 
8340=>X"00000029000000290000002900000029", 8341=>X"00000029000000290000002900000029", 8342=>X"00000028000000280000002900000029", 8343=>X"00000028000000280000002800000028", 8344=>X"00000028000000280000002800000028", 
8345=>X"00000028000000280000002800000028", 8346=>X"00000028000000280000002800000028", 8347=>X"00000028000000280000002800000028", 8348=>X"00000028000000280000002800000028", 8349=>X"00000028000000280000002800000028", 
8350=>X"00000028000000280000002800000028", 8351=>X"00000028000000280000002800000028", 8352=>X"00000028000000280000002800000028", 8353=>X"00000028000000280000002800000028", 8354=>X"00000028000000280000002800000028", 
8355=>X"00000028000000280000002800000028", 8356=>X"00000028000000280000002800000028", 8357=>X"00000028000000280000002800000028", 8358=>X"00000028000000280000002800000028", 8359=>X"00000028000000280000002800000028", 
8360=>X"00000028000000280000002800000028", 8361=>X"00000028000000280000002800000028", 8362=>X"00000028000000280000002800000028", 8363=>X"00000028000000280000002800000028", 8364=>X"00000028000000280000002800000028", 
8365=>X"00000028000000280000002800000028", 8366=>X"00000028000000280000002800000028", 8367=>X"00000028000000280000002800000028", 8368=>X"00000028000000280000002800000028", 8369=>X"00000028000000280000002800000028", 
8370=>X"00000028000000280000002800000028", 8371=>X"00000028000000280000002800000028", 8372=>X"00000028000000280000002800000028", 8373=>X"00000028000000280000002800000028", 8374=>X"00000028000000280000002800000028", 
8375=>X"00000028000000280000002800000028", 8376=>X"00000028000000280000002800000028", 8377=>X"00000028000000280000002800000028", 8378=>X"00000028000000280000002800000028", 8379=>X"00000028000000280000002800000028", 
8380=>X"00000028000000280000002800000028", 8381=>X"00000028000000280000002800000028", 8382=>X"00000028000000280000002800000028", 8383=>X"00000028000000280000002800000028", 8384=>X"00000028000000280000002800000028", 
8385=>X"00000028000000280000002800000028", 8386=>X"00000028000000280000002800000028", 8387=>X"00000028000000280000002800000028", 8388=>X"00000028000000280000002800000028", 8389=>X"00000028000000280000002800000028", 
8390=>X"00000028000000280000002800000028", 8391=>X"00000028000000280000002800000028", 8392=>X"00000028000000280000002800000028", 8393=>X"00000028000000280000002800000028", 8394=>X"00000028000000280000002800000028", 
8395=>X"00000028000000280000002800000028", 8396=>X"00000028000000280000002800000028", 8397=>X"00000028000000280000002800000028", 8398=>X"00000028000000280000002800000028", 8399=>X"00000028000000280000002800000028", 
8400=>X"00000028000000280000002800000028", 8401=>X"00000028000000280000002800000028", 8402=>X"00000028000000280000002800000028", 8403=>X"00000028000000280000002800000028", 8404=>X"00000028000000280000002800000028", 
8405=>X"00000028000000280000002800000028", 8406=>X"00000028000000280000002800000028", 8407=>X"00000028000000280000002800000028", 8408=>X"00000028000000280000002800000028", 8409=>X"00000028000000280000002800000028", 
8410=>X"00000028000000280000002800000028", 8411=>X"00000028000000280000002800000028", 8412=>X"00000028000000280000002800000028", 8413=>X"00000028000000280000002800000028", 8414=>X"00000028000000280000002800000028", 
8415=>X"00000028000000280000002800000028", 8416=>X"00000028000000280000002800000028", 8417=>X"00000028000000280000002800000028", 8418=>X"00000028000000280000002800000028", 8419=>X"00000028000000280000002800000028", 
8420=>X"00000028000000280000002800000028", 8421=>X"00000028000000280000002800000028", 8422=>X"00000028000000280000002800000028", 8423=>X"00000028000000280000002800000028", 8424=>X"00000028000000280000002800000028", 
8425=>X"00000028000000280000002800000028", 8426=>X"00000028000000280000002800000028", 8427=>X"00000028000000280000002800000028", 8428=>X"00000028000000280000002800000028", 8429=>X"00000028000000280000002800000028", 
8430=>X"00000028000000280000002800000028", 8431=>X"00000028000000280000002800000028", 8432=>X"00000028000000280000002800000028", 8433=>X"00000028000000280000002800000028", 8434=>X"00000028000000280000002800000028", 
8435=>X"00000028000000280000002800000028", 8436=>X"00000028000000280000002800000028", 8437=>X"00000028000000280000002800000028", 8438=>X"00000028000000280000002800000028", 8439=>X"00000028000000280000002800000028", 
8440=>X"00000028000000280000002800000028", 8441=>X"00000028000000280000002800000028", 8442=>X"00000028000000280000002800000028", 8443=>X"00000028000000280000002800000028", 8444=>X"00000028000000280000002800000028", 
8445=>X"00000028000000280000002800000028", 8446=>X"00000028000000280000002800000028", 8447=>X"00000028000000280000002800000028", 8448=>X"00000028000000280000002800000028", 8449=>X"00000028000000280000002800000028", 
8450=>X"00000028000000280000002800000028", 8451=>X"00000028000000280000002800000028", 8452=>X"00000028000000280000002800000028", 8453=>X"00000028000000280000002800000028", 8454=>X"00000028000000280000002800000028", 
8455=>X"00000028000000280000002800000028", 8456=>X"00000028000000280000002800000028", 8457=>X"00000028000000280000002800000028", 8458=>X"00000028000000280000002800000028", 8459=>X"00000028000000280000002800000028", 
8460=>X"00000028000000280000002800000028", 8461=>X"00000028000000280000002800000028", 8462=>X"00000028000000280000002800000028", 8463=>X"00000028000000280000002800000028", 8464=>X"00000028000000280000002800000028", 
8465=>X"00000028000000280000002800000028", 8466=>X"00000028000000280000002800000028", 8467=>X"00000028000000280000002800000028", 8468=>X"00000028000000280000002800000028", 8469=>X"00000028000000280000002800000028", 
8470=>X"00000028000000280000002800000028", 8471=>X"00000028000000280000002800000028", 8472=>X"00000028000000280000002800000028", 8473=>X"00000028000000280000002800000028", 8474=>X"00000028000000280000002800000028", 
8475=>X"00000028000000280000002800000028", 8476=>X"00000028000000280000002800000028", 8477=>X"00000028000000280000002800000028", 8478=>X"00000028000000280000002800000028", 8479=>X"00000028000000280000002800000028", 
8480=>X"00000028000000280000002800000028", 8481=>X"00000028000000280000002800000028", 8482=>X"00000028000000280000002800000028", 8483=>X"00000028000000280000002800000028", 8484=>X"00000028000000280000002800000028", 
8485=>X"00000028000000280000002800000028", 8486=>X"00000028000000280000002800000028", 8487=>X"00000028000000280000002800000028", 8488=>X"00000028000000280000002800000028", 8489=>X"00000028000000280000002800000028", 
8490=>X"00000028000000280000002800000028", 8491=>X"00000028000000280000002800000028", 8492=>X"00000028000000280000002800000028", 8493=>X"00000028000000280000002800000028", 8494=>X"00000028000000280000002800000028", 
8495=>X"00000028000000280000002800000028", 8496=>X"00000028000000280000002800000028", 8497=>X"00000028000000280000002800000028", 8498=>X"00000028000000280000002800000028", 8499=>X"00000028000000280000002800000028", 
8500=>X"00000028000000280000002800000028", 8501=>X"00000028000000280000002800000028", 8502=>X"00000028000000280000002800000028", 8503=>X"00000028000000280000002800000028", 8504=>X"00000028000000280000002800000028", 
8505=>X"00000028000000280000002800000028", 8506=>X"00000027000000270000002800000028", 8507=>X"00000027000000270000002700000027", 8508=>X"00000027000000270000002700000027", 8509=>X"00000027000000270000002700000027", 
8510=>X"00000027000000270000002700000027", 8511=>X"00000027000000270000002700000027", 8512=>X"00000027000000270000002700000027", 8513=>X"00000027000000270000002700000027", 8514=>X"00000027000000270000002700000027", 
8515=>X"00000027000000270000002700000027", 8516=>X"00000027000000270000002700000027", 8517=>X"00000027000000270000002700000027", 8518=>X"00000027000000270000002700000027", 8519=>X"00000027000000270000002700000027", 
8520=>X"00000027000000270000002700000027", 8521=>X"00000027000000270000002700000027", 8522=>X"00000027000000270000002700000027", 8523=>X"00000027000000270000002700000027", 8524=>X"00000027000000270000002700000027", 
8525=>X"00000027000000270000002700000027", 8526=>X"00000027000000270000002700000027", 8527=>X"00000027000000270000002700000027", 8528=>X"00000027000000270000002700000027", 8529=>X"00000027000000270000002700000027", 
8530=>X"00000027000000270000002700000027", 8531=>X"00000027000000270000002700000027", 8532=>X"00000027000000270000002700000027", 8533=>X"00000027000000270000002700000027", 8534=>X"00000027000000270000002700000027", 
8535=>X"00000027000000270000002700000027", 8536=>X"00000027000000270000002700000027", 8537=>X"00000027000000270000002700000027", 8538=>X"00000027000000270000002700000027", 8539=>X"00000027000000270000002700000027", 
8540=>X"00000027000000270000002700000027", 8541=>X"00000027000000270000002700000027", 8542=>X"00000027000000270000002700000027", 8543=>X"00000027000000270000002700000027", 8544=>X"00000027000000270000002700000027", 
8545=>X"00000027000000270000002700000027", 8546=>X"00000027000000270000002700000027", 8547=>X"00000027000000270000002700000027", 8548=>X"00000027000000270000002700000027", 8549=>X"00000027000000270000002700000027", 
8550=>X"00000027000000270000002700000027", 8551=>X"00000027000000270000002700000027", 8552=>X"00000027000000270000002700000027", 8553=>X"00000027000000270000002700000027", 8554=>X"00000027000000270000002700000027", 
8555=>X"00000027000000270000002700000027", 8556=>X"00000027000000270000002700000027", 8557=>X"00000027000000270000002700000027", 8558=>X"00000027000000270000002700000027", 8559=>X"00000027000000270000002700000027", 
8560=>X"00000027000000270000002700000027", 8561=>X"00000027000000270000002700000027", 8562=>X"00000027000000270000002700000027", 8563=>X"00000027000000270000002700000027", 8564=>X"00000027000000270000002700000027", 
8565=>X"00000027000000270000002700000027", 8566=>X"00000027000000270000002700000027", 8567=>X"00000027000000270000002700000027", 8568=>X"00000027000000270000002700000027", 8569=>X"00000027000000270000002700000027", 
8570=>X"00000027000000270000002700000027", 8571=>X"00000027000000270000002700000027", 8572=>X"00000027000000270000002700000027", 8573=>X"00000027000000270000002700000027", 8574=>X"00000027000000270000002700000027", 
8575=>X"00000027000000270000002700000027", 8576=>X"00000027000000270000002700000027", 8577=>X"00000027000000270000002700000027", 8578=>X"00000027000000270000002700000027", 8579=>X"00000027000000270000002700000027", 
8580=>X"00000027000000270000002700000027", 8581=>X"00000027000000270000002700000027", 8582=>X"00000027000000270000002700000027", 8583=>X"00000027000000270000002700000027", 8584=>X"00000027000000270000002700000027", 
8585=>X"00000027000000270000002700000027", 8586=>X"00000027000000270000002700000027", 8587=>X"00000027000000270000002700000027", 8588=>X"00000027000000270000002700000027", 8589=>X"00000027000000270000002700000027", 
8590=>X"00000027000000270000002700000027", 8591=>X"00000027000000270000002700000027", 8592=>X"00000027000000270000002700000027", 8593=>X"00000027000000270000002700000027", 8594=>X"00000027000000270000002700000027", 
8595=>X"00000027000000270000002700000027", 8596=>X"00000027000000270000002700000027", 8597=>X"00000027000000270000002700000027", 8598=>X"00000027000000270000002700000027", 8599=>X"00000027000000270000002700000027", 
8600=>X"00000027000000270000002700000027", 8601=>X"00000027000000270000002700000027", 8602=>X"00000027000000270000002700000027", 8603=>X"00000027000000270000002700000027", 8604=>X"00000027000000270000002700000027", 
8605=>X"00000027000000270000002700000027", 8606=>X"00000027000000270000002700000027", 8607=>X"00000027000000270000002700000027", 8608=>X"00000027000000270000002700000027", 8609=>X"00000027000000270000002700000027", 
8610=>X"00000027000000270000002700000027", 8611=>X"00000027000000270000002700000027", 8612=>X"00000027000000270000002700000027", 8613=>X"00000027000000270000002700000027", 8614=>X"00000027000000270000002700000027", 
8615=>X"00000027000000270000002700000027", 8616=>X"00000027000000270000002700000027", 8617=>X"00000027000000270000002700000027", 8618=>X"00000027000000270000002700000027", 8619=>X"00000027000000270000002700000027", 
8620=>X"00000027000000270000002700000027", 8621=>X"00000027000000270000002700000027", 8622=>X"00000027000000270000002700000027", 8623=>X"00000027000000270000002700000027", 8624=>X"00000027000000270000002700000027", 
8625=>X"00000027000000270000002700000027", 8626=>X"00000027000000270000002700000027", 8627=>X"00000027000000270000002700000027", 8628=>X"00000027000000270000002700000027", 8629=>X"00000027000000270000002700000027", 
8630=>X"00000027000000270000002700000027", 8631=>X"00000027000000270000002700000027", 8632=>X"00000027000000270000002700000027", 8633=>X"00000027000000270000002700000027", 8634=>X"00000027000000270000002700000027", 
8635=>X"00000027000000270000002700000027", 8636=>X"00000027000000270000002700000027", 8637=>X"00000027000000270000002700000027", 8638=>X"00000027000000270000002700000027", 8639=>X"00000027000000270000002700000027", 
8640=>X"00000027000000270000002700000027", 8641=>X"00000027000000270000002700000027", 8642=>X"00000027000000270000002700000027", 8643=>X"00000027000000270000002700000027", 8644=>X"00000027000000270000002700000027", 
8645=>X"00000027000000270000002700000027", 8646=>X"00000027000000270000002700000027", 8647=>X"00000027000000270000002700000027", 8648=>X"00000027000000270000002700000027", 8649=>X"00000027000000270000002700000027", 
8650=>X"00000027000000270000002700000027", 8651=>X"00000027000000270000002700000027", 8652=>X"00000027000000270000002700000027", 8653=>X"00000027000000270000002700000027", 8654=>X"00000027000000270000002700000027", 
8655=>X"00000027000000270000002700000027", 8656=>X"00000027000000270000002700000027", 8657=>X"00000027000000270000002700000027", 8658=>X"00000027000000270000002700000027", 8659=>X"00000027000000270000002700000027", 
8660=>X"00000027000000270000002700000027", 8661=>X"00000027000000270000002700000027", 8662=>X"00000027000000270000002700000027", 8663=>X"00000027000000270000002700000027", 8664=>X"00000027000000270000002700000027", 
8665=>X"00000027000000270000002700000027", 8666=>X"00000027000000270000002700000027", 8667=>X"00000027000000270000002700000027", 8668=>X"00000027000000270000002700000027", 8669=>X"00000027000000270000002700000027", 
8670=>X"00000027000000270000002700000027", 8671=>X"00000027000000270000002700000027", 8672=>X"00000027000000270000002700000027", 8673=>X"00000027000000270000002700000027", 8674=>X"00000027000000270000002700000027", 
8675=>X"00000027000000270000002700000027", 8676=>X"00000027000000270000002700000027", 8677=>X"00000027000000270000002700000027", 8678=>X"00000026000000270000002700000027", 8679=>X"00000026000000260000002600000026", 
8680=>X"00000026000000260000002600000026", 8681=>X"00000026000000260000002600000026", 8682=>X"00000026000000260000002600000026", 8683=>X"00000026000000260000002600000026", 8684=>X"00000026000000260000002600000026", 
8685=>X"00000026000000260000002600000026", 8686=>X"00000026000000260000002600000026", 8687=>X"00000026000000260000002600000026", 8688=>X"00000026000000260000002600000026", 8689=>X"00000026000000260000002600000026", 
8690=>X"00000026000000260000002600000026", 8691=>X"00000026000000260000002600000026", 8692=>X"00000026000000260000002600000026", 8693=>X"00000026000000260000002600000026", 8694=>X"00000026000000260000002600000026", 
8695=>X"00000026000000260000002600000026", 8696=>X"00000026000000260000002600000026", 8697=>X"00000026000000260000002600000026", 8698=>X"00000026000000260000002600000026", 8699=>X"00000026000000260000002600000026", 
8700=>X"00000026000000260000002600000026", 8701=>X"00000026000000260000002600000026", 8702=>X"00000026000000260000002600000026", 8703=>X"00000026000000260000002600000026", 8704=>X"00000026000000260000002600000026", 
8705=>X"00000026000000260000002600000026", 8706=>X"00000026000000260000002600000026", 8707=>X"00000026000000260000002600000026", 8708=>X"00000026000000260000002600000026", 8709=>X"00000026000000260000002600000026", 
8710=>X"00000026000000260000002600000026", 8711=>X"00000026000000260000002600000026", 8712=>X"00000026000000260000002600000026", 8713=>X"00000026000000260000002600000026", 8714=>X"00000026000000260000002600000026", 
8715=>X"00000026000000260000002600000026", 8716=>X"00000026000000260000002600000026", 8717=>X"00000026000000260000002600000026", 8718=>X"00000026000000260000002600000026", 8719=>X"00000026000000260000002600000026", 
8720=>X"00000026000000260000002600000026", 8721=>X"00000026000000260000002600000026", 8722=>X"00000026000000260000002600000026", 8723=>X"00000026000000260000002600000026", 8724=>X"00000026000000260000002600000026", 
8725=>X"00000026000000260000002600000026", 8726=>X"00000026000000260000002600000026", 8727=>X"00000026000000260000002600000026", 8728=>X"00000026000000260000002600000026", 8729=>X"00000026000000260000002600000026", 
8730=>X"00000026000000260000002600000026", 8731=>X"00000026000000260000002600000026", 8732=>X"00000026000000260000002600000026", 8733=>X"00000026000000260000002600000026", 8734=>X"00000026000000260000002600000026", 
8735=>X"00000026000000260000002600000026", 8736=>X"00000026000000260000002600000026", 8737=>X"00000026000000260000002600000026", 8738=>X"00000026000000260000002600000026", 8739=>X"00000026000000260000002600000026", 
8740=>X"00000026000000260000002600000026", 8741=>X"00000026000000260000002600000026", 8742=>X"00000026000000260000002600000026", 8743=>X"00000026000000260000002600000026", 8744=>X"00000026000000260000002600000026", 
8745=>X"00000026000000260000002600000026", 8746=>X"00000026000000260000002600000026", 8747=>X"00000026000000260000002600000026", 8748=>X"00000026000000260000002600000026", 8749=>X"00000026000000260000002600000026", 
8750=>X"00000026000000260000002600000026", 8751=>X"00000026000000260000002600000026", 8752=>X"00000026000000260000002600000026", 8753=>X"00000026000000260000002600000026", 8754=>X"00000026000000260000002600000026", 
8755=>X"00000026000000260000002600000026", 8756=>X"00000026000000260000002600000026", 8757=>X"00000026000000260000002600000026", 8758=>X"00000026000000260000002600000026", 8759=>X"00000026000000260000002600000026", 
8760=>X"00000026000000260000002600000026", 8761=>X"00000026000000260000002600000026", 8762=>X"00000026000000260000002600000026", 8763=>X"00000026000000260000002600000026", 8764=>X"00000026000000260000002600000026", 
8765=>X"00000026000000260000002600000026", 8766=>X"00000026000000260000002600000026", 8767=>X"00000026000000260000002600000026", 8768=>X"00000026000000260000002600000026", 8769=>X"00000026000000260000002600000026", 
8770=>X"00000026000000260000002600000026", 8771=>X"00000026000000260000002600000026", 8772=>X"00000026000000260000002600000026", 8773=>X"00000026000000260000002600000026", 8774=>X"00000026000000260000002600000026", 
8775=>X"00000026000000260000002600000026", 8776=>X"00000026000000260000002600000026", 8777=>X"00000026000000260000002600000026", 8778=>X"00000026000000260000002600000026", 8779=>X"00000026000000260000002600000026", 
8780=>X"00000026000000260000002600000026", 8781=>X"00000026000000260000002600000026", 8782=>X"00000026000000260000002600000026", 8783=>X"00000026000000260000002600000026", 8784=>X"00000026000000260000002600000026", 
8785=>X"00000026000000260000002600000026", 8786=>X"00000026000000260000002600000026", 8787=>X"00000026000000260000002600000026", 8788=>X"00000026000000260000002600000026", 8789=>X"00000026000000260000002600000026", 
8790=>X"00000026000000260000002600000026", 8791=>X"00000026000000260000002600000026", 8792=>X"00000026000000260000002600000026", 8793=>X"00000026000000260000002600000026", 8794=>X"00000026000000260000002600000026", 
8795=>X"00000026000000260000002600000026", 8796=>X"00000026000000260000002600000026", 8797=>X"00000026000000260000002600000026", 8798=>X"00000026000000260000002600000026", 8799=>X"00000026000000260000002600000026", 
8800=>X"00000026000000260000002600000026", 8801=>X"00000026000000260000002600000026", 8802=>X"00000026000000260000002600000026", 8803=>X"00000026000000260000002600000026", 8804=>X"00000026000000260000002600000026", 
8805=>X"00000026000000260000002600000026", 8806=>X"00000026000000260000002600000026", 8807=>X"00000026000000260000002600000026", 8808=>X"00000026000000260000002600000026", 8809=>X"00000026000000260000002600000026", 
8810=>X"00000026000000260000002600000026", 8811=>X"00000026000000260000002600000026", 8812=>X"00000026000000260000002600000026", 8813=>X"00000026000000260000002600000026", 8814=>X"00000026000000260000002600000026", 
8815=>X"00000026000000260000002600000026", 8816=>X"00000026000000260000002600000026", 8817=>X"00000026000000260000002600000026", 8818=>X"00000026000000260000002600000026", 8819=>X"00000026000000260000002600000026", 
8820=>X"00000026000000260000002600000026", 8821=>X"00000026000000260000002600000026", 8822=>X"00000026000000260000002600000026", 8823=>X"00000026000000260000002600000026", 8824=>X"00000026000000260000002600000026", 
8825=>X"00000026000000260000002600000026", 8826=>X"00000026000000260000002600000026", 8827=>X"00000026000000260000002600000026", 8828=>X"00000026000000260000002600000026", 8829=>X"00000026000000260000002600000026", 
8830=>X"00000026000000260000002600000026", 8831=>X"00000026000000260000002600000026", 8832=>X"00000026000000260000002600000026", 8833=>X"00000026000000260000002600000026", 8834=>X"00000026000000260000002600000026", 
8835=>X"00000026000000260000002600000026", 8836=>X"00000026000000260000002600000026", 8837=>X"00000026000000260000002600000026", 8838=>X"00000026000000260000002600000026", 8839=>X"00000026000000260000002600000026", 
8840=>X"00000026000000260000002600000026", 8841=>X"00000026000000260000002600000026", 8842=>X"00000026000000260000002600000026", 8843=>X"00000026000000260000002600000026", 8844=>X"00000026000000260000002600000026", 
8845=>X"00000026000000260000002600000026", 8846=>X"00000026000000260000002600000026", 8847=>X"00000026000000260000002600000026", 8848=>X"00000026000000260000002600000026", 8849=>X"00000026000000260000002600000026", 
8850=>X"00000026000000260000002600000026", 8851=>X"00000026000000260000002600000026", 8852=>X"00000026000000260000002600000026", 8853=>X"00000026000000260000002600000026", 8854=>X"00000026000000260000002600000026", 
8855=>X"00000026000000260000002600000026", 8856=>X"00000026000000260000002600000026", 8857=>X"00000026000000260000002600000026", 8858=>X"00000026000000260000002600000026", 8859=>X"00000026000000260000002600000026", 
8860=>X"00000025000000250000002600000026", 8861=>X"00000025000000250000002500000025", 8862=>X"00000025000000250000002500000025", 8863=>X"00000025000000250000002500000025", 8864=>X"00000025000000250000002500000025", 
8865=>X"00000025000000250000002500000025", 8866=>X"00000025000000250000002500000025", 8867=>X"00000025000000250000002500000025", 8868=>X"00000025000000250000002500000025", 8869=>X"00000025000000250000002500000025", 
8870=>X"00000025000000250000002500000025", 8871=>X"00000025000000250000002500000025", 8872=>X"00000025000000250000002500000025", 8873=>X"00000025000000250000002500000025", 8874=>X"00000025000000250000002500000025", 
8875=>X"00000025000000250000002500000025", 8876=>X"00000025000000250000002500000025", 8877=>X"00000025000000250000002500000025", 8878=>X"00000025000000250000002500000025", 8879=>X"00000025000000250000002500000025", 
8880=>X"00000025000000250000002500000025", 8881=>X"00000025000000250000002500000025", 8882=>X"00000025000000250000002500000025", 8883=>X"00000025000000250000002500000025", 8884=>X"00000025000000250000002500000025", 
8885=>X"00000025000000250000002500000025", 8886=>X"00000025000000250000002500000025", 8887=>X"00000025000000250000002500000025", 8888=>X"00000025000000250000002500000025", 8889=>X"00000025000000250000002500000025", 
8890=>X"00000025000000250000002500000025", 8891=>X"00000025000000250000002500000025", 8892=>X"00000025000000250000002500000025", 8893=>X"00000025000000250000002500000025", 8894=>X"00000025000000250000002500000025", 
8895=>X"00000025000000250000002500000025", 8896=>X"00000025000000250000002500000025", 8897=>X"00000025000000250000002500000025", 8898=>X"00000025000000250000002500000025", 8899=>X"00000025000000250000002500000025", 
8900=>X"00000025000000250000002500000025", 8901=>X"00000025000000250000002500000025", 8902=>X"00000025000000250000002500000025", 8903=>X"00000025000000250000002500000025", 8904=>X"00000025000000250000002500000025", 
8905=>X"00000025000000250000002500000025", 8906=>X"00000025000000250000002500000025", 8907=>X"00000025000000250000002500000025", 8908=>X"00000025000000250000002500000025", 8909=>X"00000025000000250000002500000025", 
8910=>X"00000025000000250000002500000025", 8911=>X"00000025000000250000002500000025", 8912=>X"00000025000000250000002500000025", 8913=>X"00000025000000250000002500000025", 8914=>X"00000025000000250000002500000025", 
8915=>X"00000025000000250000002500000025", 8916=>X"00000025000000250000002500000025", 8917=>X"00000025000000250000002500000025", 8918=>X"00000025000000250000002500000025", 8919=>X"00000025000000250000002500000025", 
8920=>X"00000025000000250000002500000025", 8921=>X"00000025000000250000002500000025", 8922=>X"00000025000000250000002500000025", 8923=>X"00000025000000250000002500000025", 8924=>X"00000025000000250000002500000025", 
8925=>X"00000025000000250000002500000025", 8926=>X"00000025000000250000002500000025", 8927=>X"00000025000000250000002500000025", 8928=>X"00000025000000250000002500000025", 8929=>X"00000025000000250000002500000025", 
8930=>X"00000025000000250000002500000025", 8931=>X"00000025000000250000002500000025", 8932=>X"00000025000000250000002500000025", 8933=>X"00000025000000250000002500000025", 8934=>X"00000025000000250000002500000025", 
8935=>X"00000025000000250000002500000025", 8936=>X"00000025000000250000002500000025", 8937=>X"00000025000000250000002500000025", 8938=>X"00000025000000250000002500000025", 8939=>X"00000025000000250000002500000025", 
8940=>X"00000025000000250000002500000025", 8941=>X"00000025000000250000002500000025", 8942=>X"00000025000000250000002500000025", 8943=>X"00000025000000250000002500000025", 8944=>X"00000025000000250000002500000025", 
8945=>X"00000025000000250000002500000025", 8946=>X"00000025000000250000002500000025", 8947=>X"00000025000000250000002500000025", 8948=>X"00000025000000250000002500000025", 8949=>X"00000025000000250000002500000025", 
8950=>X"00000025000000250000002500000025", 8951=>X"00000025000000250000002500000025", 8952=>X"00000025000000250000002500000025", 8953=>X"00000025000000250000002500000025", 8954=>X"00000025000000250000002500000025", 
8955=>X"00000025000000250000002500000025", 8956=>X"00000025000000250000002500000025", 8957=>X"00000025000000250000002500000025", 8958=>X"00000025000000250000002500000025", 8959=>X"00000025000000250000002500000025", 
8960=>X"00000025000000250000002500000025", 8961=>X"00000025000000250000002500000025", 8962=>X"00000025000000250000002500000025", 8963=>X"00000025000000250000002500000025", 8964=>X"00000025000000250000002500000025", 
8965=>X"00000025000000250000002500000025", 8966=>X"00000025000000250000002500000025", 8967=>X"00000025000000250000002500000025", 8968=>X"00000025000000250000002500000025", 8969=>X"00000025000000250000002500000025", 
8970=>X"00000025000000250000002500000025", 8971=>X"00000025000000250000002500000025", 8972=>X"00000025000000250000002500000025", 8973=>X"00000025000000250000002500000025", 8974=>X"00000025000000250000002500000025", 
8975=>X"00000025000000250000002500000025", 8976=>X"00000025000000250000002500000025", 8977=>X"00000025000000250000002500000025", 8978=>X"00000025000000250000002500000025", 8979=>X"00000025000000250000002500000025", 
8980=>X"00000025000000250000002500000025", 8981=>X"00000025000000250000002500000025", 8982=>X"00000025000000250000002500000025", 8983=>X"00000025000000250000002500000025", 8984=>X"00000025000000250000002500000025", 
8985=>X"00000025000000250000002500000025", 8986=>X"00000025000000250000002500000025", 8987=>X"00000025000000250000002500000025", 8988=>X"00000025000000250000002500000025", 8989=>X"00000025000000250000002500000025", 
8990=>X"00000025000000250000002500000025", 8991=>X"00000025000000250000002500000025", 8992=>X"00000025000000250000002500000025", 8993=>X"00000025000000250000002500000025", 8994=>X"00000025000000250000002500000025", 
8995=>X"00000025000000250000002500000025", 8996=>X"00000025000000250000002500000025", 8997=>X"00000025000000250000002500000025", 8998=>X"00000025000000250000002500000025", 8999=>X"00000025000000250000002500000025", 
9000=>X"00000025000000250000002500000025", 9001=>X"00000025000000250000002500000025", 9002=>X"00000025000000250000002500000025", 9003=>X"00000025000000250000002500000025", 9004=>X"00000025000000250000002500000025", 
9005=>X"00000025000000250000002500000025", 9006=>X"00000025000000250000002500000025", 9007=>X"00000025000000250000002500000025", 9008=>X"00000025000000250000002500000025", 9009=>X"00000025000000250000002500000025", 
9010=>X"00000025000000250000002500000025", 9011=>X"00000025000000250000002500000025", 9012=>X"00000025000000250000002500000025", 9013=>X"00000025000000250000002500000025", 9014=>X"00000025000000250000002500000025", 
9015=>X"00000025000000250000002500000025", 9016=>X"00000025000000250000002500000025", 9017=>X"00000025000000250000002500000025", 9018=>X"00000025000000250000002500000025", 9019=>X"00000025000000250000002500000025", 
9020=>X"00000025000000250000002500000025", 9021=>X"00000025000000250000002500000025", 9022=>X"00000025000000250000002500000025", 9023=>X"00000025000000250000002500000025", 9024=>X"00000025000000250000002500000025", 
9025=>X"00000025000000250000002500000025", 9026=>X"00000025000000250000002500000025", 9027=>X"00000025000000250000002500000025", 9028=>X"00000025000000250000002500000025", 9029=>X"00000025000000250000002500000025", 
9030=>X"00000025000000250000002500000025", 9031=>X"00000025000000250000002500000025", 9032=>X"00000025000000250000002500000025", 9033=>X"00000025000000250000002500000025", 9034=>X"00000025000000250000002500000025", 
9035=>X"00000025000000250000002500000025", 9036=>X"00000025000000250000002500000025", 9037=>X"00000025000000250000002500000025", 9038=>X"00000025000000250000002500000025", 9039=>X"00000025000000250000002500000025", 
9040=>X"00000025000000250000002500000025", 9041=>X"00000025000000250000002500000025", 9042=>X"00000025000000250000002500000025", 9043=>X"00000025000000250000002500000025", 9044=>X"00000025000000250000002500000025", 
9045=>X"00000025000000250000002500000025", 9046=>X"00000025000000250000002500000025", 9047=>X"00000025000000250000002500000025", 9048=>X"00000025000000250000002500000025", 9049=>X"00000025000000250000002500000025", 
9050=>X"00000025000000250000002500000025", 9051=>X"00000025000000250000002500000025", 9052=>X"00000024000000240000002400000024", 9053=>X"00000024000000240000002400000024", 9054=>X"00000024000000240000002400000024", 
9055=>X"00000024000000240000002400000024", 9056=>X"00000024000000240000002400000024", 9057=>X"00000024000000240000002400000024", 9058=>X"00000024000000240000002400000024", 9059=>X"00000024000000240000002400000024", 
9060=>X"00000024000000240000002400000024", 9061=>X"00000024000000240000002400000024", 9062=>X"00000024000000240000002400000024", 9063=>X"00000024000000240000002400000024", 9064=>X"00000024000000240000002400000024", 
9065=>X"00000024000000240000002400000024", 9066=>X"00000024000000240000002400000024", 9067=>X"00000024000000240000002400000024", 9068=>X"00000024000000240000002400000024", 9069=>X"00000024000000240000002400000024", 
9070=>X"00000024000000240000002400000024", 9071=>X"00000024000000240000002400000024", 9072=>X"00000024000000240000002400000024", 9073=>X"00000024000000240000002400000024", 9074=>X"00000024000000240000002400000024", 
9075=>X"00000024000000240000002400000024", 9076=>X"00000024000000240000002400000024", 9077=>X"00000024000000240000002400000024", 9078=>X"00000024000000240000002400000024", 9079=>X"00000024000000240000002400000024", 
9080=>X"00000024000000240000002400000024", 9081=>X"00000024000000240000002400000024", 9082=>X"00000024000000240000002400000024", 9083=>X"00000024000000240000002400000024", 9084=>X"00000024000000240000002400000024", 
9085=>X"00000024000000240000002400000024", 9086=>X"00000024000000240000002400000024", 9087=>X"00000024000000240000002400000024", 9088=>X"00000024000000240000002400000024", 9089=>X"00000024000000240000002400000024", 
9090=>X"00000024000000240000002400000024", 9091=>X"00000024000000240000002400000024", 9092=>X"00000024000000240000002400000024", 9093=>X"00000024000000240000002400000024", 9094=>X"00000024000000240000002400000024", 
9095=>X"00000024000000240000002400000024", 9096=>X"00000024000000240000002400000024", 9097=>X"00000024000000240000002400000024", 9098=>X"00000024000000240000002400000024", 9099=>X"00000024000000240000002400000024", 
9100=>X"00000024000000240000002400000024", 9101=>X"00000024000000240000002400000024", 9102=>X"00000024000000240000002400000024", 9103=>X"00000024000000240000002400000024", 9104=>X"00000024000000240000002400000024", 
9105=>X"00000024000000240000002400000024", 9106=>X"00000024000000240000002400000024", 9107=>X"00000024000000240000002400000024", 9108=>X"00000024000000240000002400000024", 9109=>X"00000024000000240000002400000024", 
9110=>X"00000024000000240000002400000024", 9111=>X"00000024000000240000002400000024", 9112=>X"00000024000000240000002400000024", 9113=>X"00000024000000240000002400000024", 9114=>X"00000024000000240000002400000024", 
9115=>X"00000024000000240000002400000024", 9116=>X"00000024000000240000002400000024", 9117=>X"00000024000000240000002400000024", 9118=>X"00000024000000240000002400000024", 9119=>X"00000024000000240000002400000024", 
9120=>X"00000024000000240000002400000024", 9121=>X"00000024000000240000002400000024", 9122=>X"00000024000000240000002400000024", 9123=>X"00000024000000240000002400000024", 9124=>X"00000024000000240000002400000024", 
9125=>X"00000024000000240000002400000024", 9126=>X"00000024000000240000002400000024", 9127=>X"00000024000000240000002400000024", 9128=>X"00000024000000240000002400000024", 9129=>X"00000024000000240000002400000024", 
9130=>X"00000024000000240000002400000024", 9131=>X"00000024000000240000002400000024", 9132=>X"00000024000000240000002400000024", 9133=>X"00000024000000240000002400000024", 9134=>X"00000024000000240000002400000024", 
9135=>X"00000024000000240000002400000024", 9136=>X"00000024000000240000002400000024", 9137=>X"00000024000000240000002400000024", 9138=>X"00000024000000240000002400000024", 9139=>X"00000024000000240000002400000024", 
9140=>X"00000024000000240000002400000024", 9141=>X"00000024000000240000002400000024", 9142=>X"00000024000000240000002400000024", 9143=>X"00000024000000240000002400000024", 9144=>X"00000024000000240000002400000024", 
9145=>X"00000024000000240000002400000024", 9146=>X"00000024000000240000002400000024", 9147=>X"00000024000000240000002400000024", 9148=>X"00000024000000240000002400000024", 9149=>X"00000024000000240000002400000024", 
9150=>X"00000024000000240000002400000024", 9151=>X"00000024000000240000002400000024", 9152=>X"00000024000000240000002400000024", 9153=>X"00000024000000240000002400000024", 9154=>X"00000024000000240000002400000024", 
9155=>X"00000024000000240000002400000024", 9156=>X"00000024000000240000002400000024", 9157=>X"00000024000000240000002400000024", 9158=>X"00000024000000240000002400000024", 9159=>X"00000024000000240000002400000024", 
9160=>X"00000024000000240000002400000024", 9161=>X"00000024000000240000002400000024", 9162=>X"00000024000000240000002400000024", 9163=>X"00000024000000240000002400000024", 9164=>X"00000024000000240000002400000024", 
9165=>X"00000024000000240000002400000024", 9166=>X"00000024000000240000002400000024", 9167=>X"00000024000000240000002400000024", 9168=>X"00000024000000240000002400000024", 9169=>X"00000024000000240000002400000024", 
9170=>X"00000024000000240000002400000024", 9171=>X"00000024000000240000002400000024", 9172=>X"00000024000000240000002400000024", 9173=>X"00000024000000240000002400000024", 9174=>X"00000024000000240000002400000024", 
9175=>X"00000024000000240000002400000024", 9176=>X"00000024000000240000002400000024", 9177=>X"00000024000000240000002400000024", 9178=>X"00000024000000240000002400000024", 9179=>X"00000024000000240000002400000024", 
9180=>X"00000024000000240000002400000024", 9181=>X"00000024000000240000002400000024", 9182=>X"00000024000000240000002400000024", 9183=>X"00000024000000240000002400000024", 9184=>X"00000024000000240000002400000024", 
9185=>X"00000024000000240000002400000024", 9186=>X"00000024000000240000002400000024", 9187=>X"00000024000000240000002400000024", 9188=>X"00000024000000240000002400000024", 9189=>X"00000024000000240000002400000024", 
9190=>X"00000024000000240000002400000024", 9191=>X"00000024000000240000002400000024", 9192=>X"00000024000000240000002400000024", 9193=>X"00000024000000240000002400000024", 9194=>X"00000024000000240000002400000024", 
9195=>X"00000024000000240000002400000024", 9196=>X"00000024000000240000002400000024", 9197=>X"00000024000000240000002400000024", 9198=>X"00000024000000240000002400000024", 9199=>X"00000024000000240000002400000024", 
9200=>X"00000024000000240000002400000024", 9201=>X"00000024000000240000002400000024", 9202=>X"00000024000000240000002400000024", 9203=>X"00000024000000240000002400000024", 9204=>X"00000024000000240000002400000024", 
9205=>X"00000024000000240000002400000024", 9206=>X"00000024000000240000002400000024", 9207=>X"00000024000000240000002400000024", 9208=>X"00000024000000240000002400000024", 9209=>X"00000024000000240000002400000024", 
9210=>X"00000024000000240000002400000024", 9211=>X"00000024000000240000002400000024", 9212=>X"00000024000000240000002400000024", 9213=>X"00000024000000240000002400000024", 9214=>X"00000024000000240000002400000024", 
9215=>X"00000024000000240000002400000024", 9216=>X"00000024000000240000002400000024", 9217=>X"00000024000000240000002400000024", 9218=>X"00000024000000240000002400000024", 9219=>X"00000024000000240000002400000024", 
9220=>X"00000024000000240000002400000024", 9221=>X"00000024000000240000002400000024", 9222=>X"00000024000000240000002400000024", 9223=>X"00000024000000240000002400000024", 9224=>X"00000024000000240000002400000024", 
9225=>X"00000024000000240000002400000024", 9226=>X"00000024000000240000002400000024", 9227=>X"00000024000000240000002400000024", 9228=>X"00000024000000240000002400000024", 9229=>X"00000024000000240000002400000024", 
9230=>X"00000024000000240000002400000024", 9231=>X"00000024000000240000002400000024", 9232=>X"00000024000000240000002400000024", 9233=>X"00000024000000240000002400000024", 9234=>X"00000024000000240000002400000024", 
9235=>X"00000024000000240000002400000024", 9236=>X"00000024000000240000002400000024", 9237=>X"00000024000000240000002400000024", 9238=>X"00000024000000240000002400000024", 9239=>X"00000024000000240000002400000024", 
9240=>X"00000024000000240000002400000024", 9241=>X"00000024000000240000002400000024", 9242=>X"00000024000000240000002400000024", 9243=>X"00000024000000240000002400000024", 9244=>X"00000024000000240000002400000024", 
9245=>X"00000024000000240000002400000024", 9246=>X"00000024000000240000002400000024", 9247=>X"00000024000000240000002400000024", 9248=>X"00000024000000240000002400000024", 9249=>X"00000024000000240000002400000024", 
9250=>X"00000024000000240000002400000024", 9251=>X"00000024000000240000002400000024", 9252=>X"00000024000000240000002400000024", 9253=>X"00000024000000240000002400000024", 9254=>X"00000023000000230000002300000024", 
9255=>X"00000023000000230000002300000023", 9256=>X"00000023000000230000002300000023", 9257=>X"00000023000000230000002300000023", 9258=>X"00000023000000230000002300000023", 9259=>X"00000023000000230000002300000023", 
9260=>X"00000023000000230000002300000023", 9261=>X"00000023000000230000002300000023", 9262=>X"00000023000000230000002300000023", 9263=>X"00000023000000230000002300000023", 9264=>X"00000023000000230000002300000023", 
9265=>X"00000023000000230000002300000023", 9266=>X"00000023000000230000002300000023", 9267=>X"00000023000000230000002300000023", 9268=>X"00000023000000230000002300000023", 9269=>X"00000023000000230000002300000023", 
9270=>X"00000023000000230000002300000023", 9271=>X"00000023000000230000002300000023", 9272=>X"00000023000000230000002300000023", 9273=>X"00000023000000230000002300000023", 9274=>X"00000023000000230000002300000023", 
9275=>X"00000023000000230000002300000023", 9276=>X"00000023000000230000002300000023", 9277=>X"00000023000000230000002300000023", 9278=>X"00000023000000230000002300000023", 9279=>X"00000023000000230000002300000023", 
9280=>X"00000023000000230000002300000023", 9281=>X"00000023000000230000002300000023", 9282=>X"00000023000000230000002300000023", 9283=>X"00000023000000230000002300000023", 9284=>X"00000023000000230000002300000023", 
9285=>X"00000023000000230000002300000023", 9286=>X"00000023000000230000002300000023", 9287=>X"00000023000000230000002300000023", 9288=>X"00000023000000230000002300000023", 9289=>X"00000023000000230000002300000023", 
9290=>X"00000023000000230000002300000023", 9291=>X"00000023000000230000002300000023", 9292=>X"00000023000000230000002300000023", 9293=>X"00000023000000230000002300000023", 9294=>X"00000023000000230000002300000023", 
9295=>X"00000023000000230000002300000023", 9296=>X"00000023000000230000002300000023", 9297=>X"00000023000000230000002300000023", 9298=>X"00000023000000230000002300000023", 9299=>X"00000023000000230000002300000023", 
9300=>X"00000023000000230000002300000023", 9301=>X"00000023000000230000002300000023", 9302=>X"00000023000000230000002300000023", 9303=>X"00000023000000230000002300000023", 9304=>X"00000023000000230000002300000023", 
9305=>X"00000023000000230000002300000023", 9306=>X"00000023000000230000002300000023", 9307=>X"00000023000000230000002300000023", 9308=>X"00000023000000230000002300000023", 9309=>X"00000023000000230000002300000023", 
9310=>X"00000023000000230000002300000023", 9311=>X"00000023000000230000002300000023", 9312=>X"00000023000000230000002300000023", 9313=>X"00000023000000230000002300000023", 9314=>X"00000023000000230000002300000023", 
9315=>X"00000023000000230000002300000023", 9316=>X"00000023000000230000002300000023", 9317=>X"00000023000000230000002300000023", 9318=>X"00000023000000230000002300000023", 9319=>X"00000023000000230000002300000023", 
9320=>X"00000023000000230000002300000023", 9321=>X"00000023000000230000002300000023", 9322=>X"00000023000000230000002300000023", 9323=>X"00000023000000230000002300000023", 9324=>X"00000023000000230000002300000023", 
9325=>X"00000023000000230000002300000023", 9326=>X"00000023000000230000002300000023", 9327=>X"00000023000000230000002300000023", 9328=>X"00000023000000230000002300000023", 9329=>X"00000023000000230000002300000023", 
9330=>X"00000023000000230000002300000023", 9331=>X"00000023000000230000002300000023", 9332=>X"00000023000000230000002300000023", 9333=>X"00000023000000230000002300000023", 9334=>X"00000023000000230000002300000023", 
9335=>X"00000023000000230000002300000023", 9336=>X"00000023000000230000002300000023", 9337=>X"00000023000000230000002300000023", 9338=>X"00000023000000230000002300000023", 9339=>X"00000023000000230000002300000023", 
9340=>X"00000023000000230000002300000023", 9341=>X"00000023000000230000002300000023", 9342=>X"00000023000000230000002300000023", 9343=>X"00000023000000230000002300000023", 9344=>X"00000023000000230000002300000023", 
9345=>X"00000023000000230000002300000023", 9346=>X"00000023000000230000002300000023", 9347=>X"00000023000000230000002300000023", 9348=>X"00000023000000230000002300000023", 9349=>X"00000023000000230000002300000023", 
9350=>X"00000023000000230000002300000023", 9351=>X"00000023000000230000002300000023", 9352=>X"00000023000000230000002300000023", 9353=>X"00000023000000230000002300000023", 9354=>X"00000023000000230000002300000023", 
9355=>X"00000023000000230000002300000023", 9356=>X"00000023000000230000002300000023", 9357=>X"00000023000000230000002300000023", 9358=>X"00000023000000230000002300000023", 9359=>X"00000023000000230000002300000023", 
9360=>X"00000023000000230000002300000023", 9361=>X"00000023000000230000002300000023", 9362=>X"00000023000000230000002300000023", 9363=>X"00000023000000230000002300000023", 9364=>X"00000023000000230000002300000023", 
9365=>X"00000023000000230000002300000023", 9366=>X"00000023000000230000002300000023", 9367=>X"00000023000000230000002300000023", 9368=>X"00000023000000230000002300000023", 9369=>X"00000023000000230000002300000023", 
9370=>X"00000023000000230000002300000023", 9371=>X"00000023000000230000002300000023", 9372=>X"00000023000000230000002300000023", 9373=>X"00000023000000230000002300000023", 9374=>X"00000023000000230000002300000023", 
9375=>X"00000023000000230000002300000023", 9376=>X"00000023000000230000002300000023", 9377=>X"00000023000000230000002300000023", 9378=>X"00000023000000230000002300000023", 9379=>X"00000023000000230000002300000023", 
9380=>X"00000023000000230000002300000023", 9381=>X"00000023000000230000002300000023", 9382=>X"00000023000000230000002300000023", 9383=>X"00000023000000230000002300000023", 9384=>X"00000023000000230000002300000023", 
9385=>X"00000023000000230000002300000023", 9386=>X"00000023000000230000002300000023", 9387=>X"00000023000000230000002300000023", 9388=>X"00000023000000230000002300000023", 9389=>X"00000023000000230000002300000023", 
9390=>X"00000023000000230000002300000023", 9391=>X"00000023000000230000002300000023", 9392=>X"00000023000000230000002300000023", 9393=>X"00000023000000230000002300000023", 9394=>X"00000023000000230000002300000023", 
9395=>X"00000023000000230000002300000023", 9396=>X"00000023000000230000002300000023", 9397=>X"00000023000000230000002300000023", 9398=>X"00000023000000230000002300000023", 9399=>X"00000023000000230000002300000023", 
9400=>X"00000023000000230000002300000023", 9401=>X"00000023000000230000002300000023", 9402=>X"00000023000000230000002300000023", 9403=>X"00000023000000230000002300000023", 9404=>X"00000023000000230000002300000023", 
9405=>X"00000023000000230000002300000023", 9406=>X"00000023000000230000002300000023", 9407=>X"00000023000000230000002300000023", 9408=>X"00000023000000230000002300000023", 9409=>X"00000023000000230000002300000023", 
9410=>X"00000023000000230000002300000023", 9411=>X"00000023000000230000002300000023", 9412=>X"00000023000000230000002300000023", 9413=>X"00000023000000230000002300000023", 9414=>X"00000023000000230000002300000023", 
9415=>X"00000023000000230000002300000023", 9416=>X"00000023000000230000002300000023", 9417=>X"00000023000000230000002300000023", 9418=>X"00000023000000230000002300000023", 9419=>X"00000023000000230000002300000023", 
9420=>X"00000023000000230000002300000023", 9421=>X"00000023000000230000002300000023", 9422=>X"00000023000000230000002300000023", 9423=>X"00000023000000230000002300000023", 9424=>X"00000023000000230000002300000023", 
9425=>X"00000023000000230000002300000023", 9426=>X"00000023000000230000002300000023", 9427=>X"00000023000000230000002300000023", 9428=>X"00000023000000230000002300000023", 9429=>X"00000023000000230000002300000023", 
9430=>X"00000023000000230000002300000023", 9431=>X"00000023000000230000002300000023", 9432=>X"00000023000000230000002300000023", 9433=>X"00000023000000230000002300000023", 9434=>X"00000023000000230000002300000023", 
9435=>X"00000023000000230000002300000023", 9436=>X"00000023000000230000002300000023", 9437=>X"00000023000000230000002300000023", 9438=>X"00000023000000230000002300000023", 9439=>X"00000023000000230000002300000023", 
9440=>X"00000023000000230000002300000023", 9441=>X"00000023000000230000002300000023", 9442=>X"00000023000000230000002300000023", 9443=>X"00000023000000230000002300000023", 9444=>X"00000023000000230000002300000023", 
9445=>X"00000023000000230000002300000023", 9446=>X"00000023000000230000002300000023", 9447=>X"00000023000000230000002300000023", 9448=>X"00000023000000230000002300000023", 9449=>X"00000023000000230000002300000023", 
9450=>X"00000023000000230000002300000023", 9451=>X"00000023000000230000002300000023", 9452=>X"00000023000000230000002300000023", 9453=>X"00000023000000230000002300000023", 9454=>X"00000023000000230000002300000023", 
9455=>X"00000023000000230000002300000023", 9456=>X"00000023000000230000002300000023", 9457=>X"00000023000000230000002300000023", 9458=>X"00000023000000230000002300000023", 9459=>X"00000023000000230000002300000023", 
9460=>X"00000023000000230000002300000023", 9461=>X"00000023000000230000002300000023", 9462=>X"00000023000000230000002300000023", 9463=>X"00000023000000230000002300000023", 9464=>X"00000023000000230000002300000023", 
9465=>X"00000023000000230000002300000023", 9466=>X"00000023000000230000002300000023", 9467=>X"00000023000000230000002300000023", 9468=>X"00000022000000220000002200000023", 9469=>X"00000022000000220000002200000022", 
9470=>X"00000022000000220000002200000022", 9471=>X"00000022000000220000002200000022", 9472=>X"00000022000000220000002200000022", 9473=>X"00000022000000220000002200000022", 9474=>X"00000022000000220000002200000022", 
9475=>X"00000022000000220000002200000022", 9476=>X"00000022000000220000002200000022", 9477=>X"00000022000000220000002200000022", 9478=>X"00000022000000220000002200000022", 9479=>X"00000022000000220000002200000022", 
9480=>X"00000022000000220000002200000022", 9481=>X"00000022000000220000002200000022", 9482=>X"00000022000000220000002200000022", 9483=>X"00000022000000220000002200000022", 9484=>X"00000022000000220000002200000022", 
9485=>X"00000022000000220000002200000022", 9486=>X"00000022000000220000002200000022", 9487=>X"00000022000000220000002200000022", 9488=>X"00000022000000220000002200000022", 9489=>X"00000022000000220000002200000022", 
9490=>X"00000022000000220000002200000022", 9491=>X"00000022000000220000002200000022", 9492=>X"00000022000000220000002200000022", 9493=>X"00000022000000220000002200000022", 9494=>X"00000022000000220000002200000022", 
9495=>X"00000022000000220000002200000022", 9496=>X"00000022000000220000002200000022", 9497=>X"00000022000000220000002200000022", 9498=>X"00000022000000220000002200000022", 9499=>X"00000022000000220000002200000022", 
9500=>X"00000022000000220000002200000022", 9501=>X"00000022000000220000002200000022", 9502=>X"00000022000000220000002200000022", 9503=>X"00000022000000220000002200000022", 9504=>X"00000022000000220000002200000022", 
9505=>X"00000022000000220000002200000022", 9506=>X"00000022000000220000002200000022", 9507=>X"00000022000000220000002200000022", 9508=>X"00000022000000220000002200000022", 9509=>X"00000022000000220000002200000022", 
9510=>X"00000022000000220000002200000022", 9511=>X"00000022000000220000002200000022", 9512=>X"00000022000000220000002200000022", 9513=>X"00000022000000220000002200000022", 9514=>X"00000022000000220000002200000022", 
9515=>X"00000022000000220000002200000022", 9516=>X"00000022000000220000002200000022", 9517=>X"00000022000000220000002200000022", 9518=>X"00000022000000220000002200000022", 9519=>X"00000022000000220000002200000022", 
9520=>X"00000022000000220000002200000022", 9521=>X"00000022000000220000002200000022", 9522=>X"00000022000000220000002200000022", 9523=>X"00000022000000220000002200000022", 9524=>X"00000022000000220000002200000022", 
9525=>X"00000022000000220000002200000022", 9526=>X"00000022000000220000002200000022", 9527=>X"00000022000000220000002200000022", 9528=>X"00000022000000220000002200000022", 9529=>X"00000022000000220000002200000022", 
9530=>X"00000022000000220000002200000022", 9531=>X"00000022000000220000002200000022", 9532=>X"00000022000000220000002200000022", 9533=>X"00000022000000220000002200000022", 9534=>X"00000022000000220000002200000022", 
9535=>X"00000022000000220000002200000022", 9536=>X"00000022000000220000002200000022", 9537=>X"00000022000000220000002200000022", 9538=>X"00000022000000220000002200000022", 9539=>X"00000022000000220000002200000022", 
9540=>X"00000022000000220000002200000022", 9541=>X"00000022000000220000002200000022", 9542=>X"00000022000000220000002200000022", 9543=>X"00000022000000220000002200000022", 9544=>X"00000022000000220000002200000022", 
9545=>X"00000022000000220000002200000022", 9546=>X"00000022000000220000002200000022", 9547=>X"00000022000000220000002200000022", 9548=>X"00000022000000220000002200000022", 9549=>X"00000022000000220000002200000022", 
9550=>X"00000022000000220000002200000022", 9551=>X"00000022000000220000002200000022", 9552=>X"00000022000000220000002200000022", 9553=>X"00000022000000220000002200000022", 9554=>X"00000022000000220000002200000022", 
9555=>X"00000022000000220000002200000022", 9556=>X"00000022000000220000002200000022", 9557=>X"00000022000000220000002200000022", 9558=>X"00000022000000220000002200000022", 9559=>X"00000022000000220000002200000022", 
9560=>X"00000022000000220000002200000022", 9561=>X"00000022000000220000002200000022", 9562=>X"00000022000000220000002200000022", 9563=>X"00000022000000220000002200000022", 9564=>X"00000022000000220000002200000022", 
9565=>X"00000022000000220000002200000022", 9566=>X"00000022000000220000002200000022", 9567=>X"00000022000000220000002200000022", 9568=>X"00000022000000220000002200000022", 9569=>X"00000022000000220000002200000022", 
9570=>X"00000022000000220000002200000022", 9571=>X"00000022000000220000002200000022", 9572=>X"00000022000000220000002200000022", 9573=>X"00000022000000220000002200000022", 9574=>X"00000022000000220000002200000022", 
9575=>X"00000022000000220000002200000022", 9576=>X"00000022000000220000002200000022", 9577=>X"00000022000000220000002200000022", 9578=>X"00000022000000220000002200000022", 9579=>X"00000022000000220000002200000022", 
9580=>X"00000022000000220000002200000022", 9581=>X"00000022000000220000002200000022", 9582=>X"00000022000000220000002200000022", 9583=>X"00000022000000220000002200000022", 9584=>X"00000022000000220000002200000022", 
9585=>X"00000022000000220000002200000022", 9586=>X"00000022000000220000002200000022", 9587=>X"00000022000000220000002200000022", 9588=>X"00000022000000220000002200000022", 9589=>X"00000022000000220000002200000022", 
9590=>X"00000022000000220000002200000022", 9591=>X"00000022000000220000002200000022", 9592=>X"00000022000000220000002200000022", 9593=>X"00000022000000220000002200000022", 9594=>X"00000022000000220000002200000022", 
9595=>X"00000022000000220000002200000022", 9596=>X"00000022000000220000002200000022", 9597=>X"00000022000000220000002200000022", 9598=>X"00000022000000220000002200000022", 9599=>X"00000022000000220000002200000022", 
9600=>X"00000022000000220000002200000022", 9601=>X"00000022000000220000002200000022", 9602=>X"00000022000000220000002200000022", 9603=>X"00000022000000220000002200000022", 9604=>X"00000022000000220000002200000022", 
9605=>X"00000022000000220000002200000022", 9606=>X"00000022000000220000002200000022", 9607=>X"00000022000000220000002200000022", 9608=>X"00000022000000220000002200000022", 9609=>X"00000022000000220000002200000022", 
9610=>X"00000022000000220000002200000022", 9611=>X"00000022000000220000002200000022", 9612=>X"00000022000000220000002200000022", 9613=>X"00000022000000220000002200000022", 9614=>X"00000022000000220000002200000022", 
9615=>X"00000022000000220000002200000022", 9616=>X"00000022000000220000002200000022", 9617=>X"00000022000000220000002200000022", 9618=>X"00000022000000220000002200000022", 9619=>X"00000022000000220000002200000022", 
9620=>X"00000022000000220000002200000022", 9621=>X"00000022000000220000002200000022", 9622=>X"00000022000000220000002200000022", 9623=>X"00000022000000220000002200000022", 9624=>X"00000022000000220000002200000022", 
9625=>X"00000022000000220000002200000022", 9626=>X"00000022000000220000002200000022", 9627=>X"00000022000000220000002200000022", 9628=>X"00000022000000220000002200000022", 9629=>X"00000022000000220000002200000022", 
9630=>X"00000022000000220000002200000022", 9631=>X"00000022000000220000002200000022", 9632=>X"00000022000000220000002200000022", 9633=>X"00000022000000220000002200000022", 9634=>X"00000022000000220000002200000022", 
9635=>X"00000022000000220000002200000022", 9636=>X"00000022000000220000002200000022", 9637=>X"00000022000000220000002200000022", 9638=>X"00000022000000220000002200000022", 9639=>X"00000022000000220000002200000022", 
9640=>X"00000022000000220000002200000022", 9641=>X"00000022000000220000002200000022", 9642=>X"00000022000000220000002200000022", 9643=>X"00000022000000220000002200000022", 9644=>X"00000022000000220000002200000022", 
9645=>X"00000022000000220000002200000022", 9646=>X"00000022000000220000002200000022", 9647=>X"00000022000000220000002200000022", 9648=>X"00000022000000220000002200000022", 9649=>X"00000022000000220000002200000022", 
9650=>X"00000022000000220000002200000022", 9651=>X"00000022000000220000002200000022", 9652=>X"00000022000000220000002200000022", 9653=>X"00000022000000220000002200000022", 9654=>X"00000022000000220000002200000022", 
9655=>X"00000022000000220000002200000022", 9656=>X"00000022000000220000002200000022", 9657=>X"00000022000000220000002200000022", 9658=>X"00000022000000220000002200000022", 9659=>X"00000022000000220000002200000022", 
9660=>X"00000022000000220000002200000022", 9661=>X"00000022000000220000002200000022", 9662=>X"00000022000000220000002200000022", 9663=>X"00000022000000220000002200000022", 9664=>X"00000022000000220000002200000022", 
9665=>X"00000022000000220000002200000022", 9666=>X"00000022000000220000002200000022", 9667=>X"00000022000000220000002200000022", 9668=>X"00000022000000220000002200000022", 9669=>X"00000022000000220000002200000022", 
9670=>X"00000022000000220000002200000022", 9671=>X"00000022000000220000002200000022", 9672=>X"00000022000000220000002200000022", 9673=>X"00000022000000220000002200000022", 9674=>X"00000022000000220000002200000022", 
9675=>X"00000022000000220000002200000022", 9676=>X"00000022000000220000002200000022", 9677=>X"00000022000000220000002200000022", 9678=>X"00000022000000220000002200000022", 9679=>X"00000022000000220000002200000022", 
9680=>X"00000022000000220000002200000022", 9681=>X"00000022000000220000002200000022", 9682=>X"00000022000000220000002200000022", 9683=>X"00000022000000220000002200000022", 9684=>X"00000022000000220000002200000022", 
9685=>X"00000022000000220000002200000022", 9686=>X"00000022000000220000002200000022", 9687=>X"00000022000000220000002200000022", 9688=>X"00000022000000220000002200000022", 9689=>X"00000022000000220000002200000022", 
9690=>X"00000022000000220000002200000022", 9691=>X"00000022000000220000002200000022", 9692=>X"00000022000000220000002200000022", 9693=>X"00000022000000220000002200000022", 9694=>X"00000022000000220000002200000022", 
9695=>X"00000021000000210000002100000021", 9696=>X"00000021000000210000002100000021", 9697=>X"00000021000000210000002100000021", 9698=>X"00000021000000210000002100000021", 9699=>X"00000021000000210000002100000021", 
9700=>X"00000021000000210000002100000021", 9701=>X"00000021000000210000002100000021", 9702=>X"00000021000000210000002100000021", 9703=>X"00000021000000210000002100000021", 9704=>X"00000021000000210000002100000021", 
9705=>X"00000021000000210000002100000021", 9706=>X"00000021000000210000002100000021", 9707=>X"00000021000000210000002100000021", 9708=>X"00000021000000210000002100000021", 9709=>X"00000021000000210000002100000021", 
9710=>X"00000021000000210000002100000021", 9711=>X"00000021000000210000002100000021", 9712=>X"00000021000000210000002100000021", 9713=>X"00000021000000210000002100000021", 9714=>X"00000021000000210000002100000021", 
9715=>X"00000021000000210000002100000021", 9716=>X"00000021000000210000002100000021", 9717=>X"00000021000000210000002100000021", 9718=>X"00000021000000210000002100000021", 9719=>X"00000021000000210000002100000021", 
9720=>X"00000021000000210000002100000021", 9721=>X"00000021000000210000002100000021", 9722=>X"00000021000000210000002100000021", 9723=>X"00000021000000210000002100000021", 9724=>X"00000021000000210000002100000021", 
9725=>X"00000021000000210000002100000021", 9726=>X"00000021000000210000002100000021", 9727=>X"00000021000000210000002100000021", 9728=>X"00000021000000210000002100000021", 9729=>X"00000021000000210000002100000021", 
9730=>X"00000021000000210000002100000021", 9731=>X"00000021000000210000002100000021", 9732=>X"00000021000000210000002100000021", 9733=>X"00000021000000210000002100000021", 9734=>X"00000021000000210000002100000021", 
9735=>X"00000021000000210000002100000021", 9736=>X"00000021000000210000002100000021", 9737=>X"00000021000000210000002100000021", 9738=>X"00000021000000210000002100000021", 9739=>X"00000021000000210000002100000021", 
9740=>X"00000021000000210000002100000021", 9741=>X"00000021000000210000002100000021", 9742=>X"00000021000000210000002100000021", 9743=>X"00000021000000210000002100000021", 9744=>X"00000021000000210000002100000021", 
9745=>X"00000021000000210000002100000021", 9746=>X"00000021000000210000002100000021", 9747=>X"00000021000000210000002100000021", 9748=>X"00000021000000210000002100000021", 9749=>X"00000021000000210000002100000021", 
9750=>X"00000021000000210000002100000021", 9751=>X"00000021000000210000002100000021", 9752=>X"00000021000000210000002100000021", 9753=>X"00000021000000210000002100000021", 9754=>X"00000021000000210000002100000021", 
9755=>X"00000021000000210000002100000021", 9756=>X"00000021000000210000002100000021", 9757=>X"00000021000000210000002100000021", 9758=>X"00000021000000210000002100000021", 9759=>X"00000021000000210000002100000021", 
9760=>X"00000021000000210000002100000021", 9761=>X"00000021000000210000002100000021", 9762=>X"00000021000000210000002100000021", 9763=>X"00000021000000210000002100000021", 9764=>X"00000021000000210000002100000021", 
9765=>X"00000021000000210000002100000021", 9766=>X"00000021000000210000002100000021", 9767=>X"00000021000000210000002100000021", 9768=>X"00000021000000210000002100000021", 9769=>X"00000021000000210000002100000021", 
9770=>X"00000021000000210000002100000021", 9771=>X"00000021000000210000002100000021", 9772=>X"00000021000000210000002100000021", 9773=>X"00000021000000210000002100000021", 9774=>X"00000021000000210000002100000021", 
9775=>X"00000021000000210000002100000021", 9776=>X"00000021000000210000002100000021", 9777=>X"00000021000000210000002100000021", 9778=>X"00000021000000210000002100000021", 9779=>X"00000021000000210000002100000021", 
9780=>X"00000021000000210000002100000021", 9781=>X"00000021000000210000002100000021", 9782=>X"00000021000000210000002100000021", 9783=>X"00000021000000210000002100000021", 9784=>X"00000021000000210000002100000021", 
9785=>X"00000021000000210000002100000021", 9786=>X"00000021000000210000002100000021", 9787=>X"00000021000000210000002100000021", 9788=>X"00000021000000210000002100000021", 9789=>X"00000021000000210000002100000021", 
9790=>X"00000021000000210000002100000021", 9791=>X"00000021000000210000002100000021", 9792=>X"00000021000000210000002100000021", 9793=>X"00000021000000210000002100000021", 9794=>X"00000021000000210000002100000021", 
9795=>X"00000021000000210000002100000021", 9796=>X"00000021000000210000002100000021", 9797=>X"00000021000000210000002100000021", 9798=>X"00000021000000210000002100000021", 9799=>X"00000021000000210000002100000021", 
9800=>X"00000021000000210000002100000021", 9801=>X"00000021000000210000002100000021", 9802=>X"00000021000000210000002100000021", 9803=>X"00000021000000210000002100000021", 9804=>X"00000021000000210000002100000021", 
9805=>X"00000021000000210000002100000021", 9806=>X"00000021000000210000002100000021", 9807=>X"00000021000000210000002100000021", 9808=>X"00000021000000210000002100000021", 9809=>X"00000021000000210000002100000021", 
9810=>X"00000021000000210000002100000021", 9811=>X"00000021000000210000002100000021", 9812=>X"00000021000000210000002100000021", 9813=>X"00000021000000210000002100000021", 9814=>X"00000021000000210000002100000021", 
9815=>X"00000021000000210000002100000021", 9816=>X"00000021000000210000002100000021", 9817=>X"00000021000000210000002100000021", 9818=>X"00000021000000210000002100000021", 9819=>X"00000021000000210000002100000021", 
9820=>X"00000021000000210000002100000021", 9821=>X"00000021000000210000002100000021", 9822=>X"00000021000000210000002100000021", 9823=>X"00000021000000210000002100000021", 9824=>X"00000021000000210000002100000021", 
9825=>X"00000021000000210000002100000021", 9826=>X"00000021000000210000002100000021", 9827=>X"00000021000000210000002100000021", 9828=>X"00000021000000210000002100000021", 9829=>X"00000021000000210000002100000021", 
9830=>X"00000021000000210000002100000021", 9831=>X"00000021000000210000002100000021", 9832=>X"00000021000000210000002100000021", 9833=>X"00000021000000210000002100000021", 9834=>X"00000021000000210000002100000021", 
9835=>X"00000021000000210000002100000021", 9836=>X"00000021000000210000002100000021", 9837=>X"00000021000000210000002100000021", 9838=>X"00000021000000210000002100000021", 9839=>X"00000021000000210000002100000021", 
9840=>X"00000021000000210000002100000021", 9841=>X"00000021000000210000002100000021", 9842=>X"00000021000000210000002100000021", 9843=>X"00000021000000210000002100000021", 9844=>X"00000021000000210000002100000021", 
9845=>X"00000021000000210000002100000021", 9846=>X"00000021000000210000002100000021", 9847=>X"00000021000000210000002100000021", 9848=>X"00000021000000210000002100000021", 9849=>X"00000021000000210000002100000021", 
9850=>X"00000021000000210000002100000021", 9851=>X"00000021000000210000002100000021", 9852=>X"00000021000000210000002100000021", 9853=>X"00000021000000210000002100000021", 9854=>X"00000021000000210000002100000021", 
9855=>X"00000021000000210000002100000021", 9856=>X"00000021000000210000002100000021", 9857=>X"00000021000000210000002100000021", 9858=>X"00000021000000210000002100000021", 9859=>X"00000021000000210000002100000021", 
9860=>X"00000021000000210000002100000021", 9861=>X"00000021000000210000002100000021", 9862=>X"00000021000000210000002100000021", 9863=>X"00000021000000210000002100000021", 9864=>X"00000021000000210000002100000021", 
9865=>X"00000021000000210000002100000021", 9866=>X"00000021000000210000002100000021", 9867=>X"00000021000000210000002100000021", 9868=>X"00000021000000210000002100000021", 9869=>X"00000021000000210000002100000021", 
9870=>X"00000021000000210000002100000021", 9871=>X"00000021000000210000002100000021", 9872=>X"00000021000000210000002100000021", 9873=>X"00000021000000210000002100000021", 9874=>X"00000021000000210000002100000021", 
9875=>X"00000021000000210000002100000021", 9876=>X"00000021000000210000002100000021", 9877=>X"00000021000000210000002100000021", 9878=>X"00000021000000210000002100000021", 9879=>X"00000021000000210000002100000021", 
9880=>X"00000021000000210000002100000021", 9881=>X"00000021000000210000002100000021", 9882=>X"00000021000000210000002100000021", 9883=>X"00000021000000210000002100000021", 9884=>X"00000021000000210000002100000021", 
9885=>X"00000021000000210000002100000021", 9886=>X"00000021000000210000002100000021", 9887=>X"00000021000000210000002100000021", 9888=>X"00000021000000210000002100000021", 9889=>X"00000021000000210000002100000021", 
9890=>X"00000021000000210000002100000021", 9891=>X"00000021000000210000002100000021", 9892=>X"00000021000000210000002100000021", 9893=>X"00000021000000210000002100000021", 9894=>X"00000021000000210000002100000021", 
9895=>X"00000021000000210000002100000021", 9896=>X"00000021000000210000002100000021", 9897=>X"00000021000000210000002100000021", 9898=>X"00000021000000210000002100000021", 9899=>X"00000021000000210000002100000021", 
9900=>X"00000021000000210000002100000021", 9901=>X"00000021000000210000002100000021", 9902=>X"00000021000000210000002100000021", 9903=>X"00000021000000210000002100000021", 9904=>X"00000021000000210000002100000021", 
9905=>X"00000021000000210000002100000021", 9906=>X"00000021000000210000002100000021", 9907=>X"00000021000000210000002100000021", 9908=>X"00000021000000210000002100000021", 9909=>X"00000021000000210000002100000021", 
9910=>X"00000021000000210000002100000021", 9911=>X"00000021000000210000002100000021", 9912=>X"00000021000000210000002100000021", 9913=>X"00000021000000210000002100000021", 9914=>X"00000021000000210000002100000021", 
9915=>X"00000021000000210000002100000021", 9916=>X"00000021000000210000002100000021", 9917=>X"00000021000000210000002100000021", 9918=>X"00000021000000210000002100000021", 9919=>X"00000021000000210000002100000021", 
9920=>X"00000021000000210000002100000021", 9921=>X"00000021000000210000002100000021", 9922=>X"00000021000000210000002100000021", 9923=>X"00000021000000210000002100000021", 9924=>X"00000021000000210000002100000021", 
9925=>X"00000021000000210000002100000021", 9926=>X"00000021000000210000002100000021", 9927=>X"00000021000000210000002100000021", 9928=>X"00000021000000210000002100000021", 9929=>X"00000021000000210000002100000021", 
9930=>X"00000021000000210000002100000021", 9931=>X"00000021000000210000002100000021", 9932=>X"00000021000000210000002100000021", 9933=>X"00000021000000210000002100000021", 9934=>X"00000021000000210000002100000021", 
9935=>X"00000020000000210000002100000021", 9936=>X"00000020000000200000002000000020", 9937=>X"00000020000000200000002000000020", 9938=>X"00000020000000200000002000000020", 9939=>X"00000020000000200000002000000020", 
9940=>X"00000020000000200000002000000020", 9941=>X"00000020000000200000002000000020", 9942=>X"00000020000000200000002000000020", 9943=>X"00000020000000200000002000000020", 9944=>X"00000020000000200000002000000020", 
9945=>X"00000020000000200000002000000020", 9946=>X"00000020000000200000002000000020", 9947=>X"00000020000000200000002000000020", 9948=>X"00000020000000200000002000000020", 9949=>X"00000020000000200000002000000020", 
9950=>X"00000020000000200000002000000020", 9951=>X"00000020000000200000002000000020", 9952=>X"00000020000000200000002000000020", 9953=>X"00000020000000200000002000000020", 9954=>X"00000020000000200000002000000020", 
9955=>X"00000020000000200000002000000020", 9956=>X"00000020000000200000002000000020", 9957=>X"00000020000000200000002000000020", 9958=>X"00000020000000200000002000000020", 9959=>X"00000020000000200000002000000020", 
9960=>X"00000020000000200000002000000020", 9961=>X"00000020000000200000002000000020", 9962=>X"00000020000000200000002000000020", 9963=>X"00000020000000200000002000000020", 9964=>X"00000020000000200000002000000020", 
9965=>X"00000020000000200000002000000020", 9966=>X"00000020000000200000002000000020", 9967=>X"00000020000000200000002000000020", 9968=>X"00000020000000200000002000000020", 9969=>X"00000020000000200000002000000020", 
9970=>X"00000020000000200000002000000020", 9971=>X"00000020000000200000002000000020", 9972=>X"00000020000000200000002000000020", 9973=>X"00000020000000200000002000000020", 9974=>X"00000020000000200000002000000020", 
9975=>X"00000020000000200000002000000020", 9976=>X"00000020000000200000002000000020", 9977=>X"00000020000000200000002000000020", 9978=>X"00000020000000200000002000000020", 9979=>X"00000020000000200000002000000020", 
9980=>X"00000020000000200000002000000020", 9981=>X"00000020000000200000002000000020", 9982=>X"00000020000000200000002000000020", 9983=>X"00000020000000200000002000000020", 9984=>X"00000020000000200000002000000020", 
9985=>X"00000020000000200000002000000020", 9986=>X"00000020000000200000002000000020", 9987=>X"00000020000000200000002000000020", 9988=>X"00000020000000200000002000000020", 9989=>X"00000020000000200000002000000020", 
9990=>X"00000020000000200000002000000020", 9991=>X"00000020000000200000002000000020", 9992=>X"00000020000000200000002000000020", 9993=>X"00000020000000200000002000000020", 9994=>X"00000020000000200000002000000020", 
9995=>X"00000020000000200000002000000020", 9996=>X"00000020000000200000002000000020", 9997=>X"00000020000000200000002000000020", 9998=>X"00000020000000200000002000000020", 9999=>X"00000020000000200000002000000020", 
10000=>X"00000020000000200000002000000020", 10001=>X"00000020000000200000002000000020", 10002=>X"00000020000000200000002000000020", 10003=>X"00000020000000200000002000000020", 10004=>X"00000020000000200000002000000020", 
10005=>X"00000020000000200000002000000020", 10006=>X"00000020000000200000002000000020", 10007=>X"00000020000000200000002000000020", 10008=>X"00000020000000200000002000000020", 10009=>X"00000020000000200000002000000020", 
10010=>X"00000020000000200000002000000020", 10011=>X"00000020000000200000002000000020", 10012=>X"00000020000000200000002000000020", 10013=>X"00000020000000200000002000000020", 10014=>X"00000020000000200000002000000020", 
10015=>X"00000020000000200000002000000020", 10016=>X"00000020000000200000002000000020", 10017=>X"00000020000000200000002000000020", 10018=>X"00000020000000200000002000000020", 10019=>X"00000020000000200000002000000020", 
10020=>X"00000020000000200000002000000020", 10021=>X"00000020000000200000002000000020", 10022=>X"00000020000000200000002000000020", 10023=>X"00000020000000200000002000000020", 10024=>X"00000020000000200000002000000020", 
10025=>X"00000020000000200000002000000020", 10026=>X"00000020000000200000002000000020", 10027=>X"00000020000000200000002000000020", 10028=>X"00000020000000200000002000000020", 10029=>X"00000020000000200000002000000020", 
10030=>X"00000020000000200000002000000020", 10031=>X"00000020000000200000002000000020", 10032=>X"00000020000000200000002000000020", 10033=>X"00000020000000200000002000000020", 10034=>X"00000020000000200000002000000020", 
10035=>X"00000020000000200000002000000020", 10036=>X"00000020000000200000002000000020", 10037=>X"00000020000000200000002000000020", 10038=>X"00000020000000200000002000000020", 10039=>X"00000020000000200000002000000020", 
10040=>X"00000020000000200000002000000020", 10041=>X"00000020000000200000002000000020", 10042=>X"00000020000000200000002000000020", 10043=>X"00000020000000200000002000000020", 10044=>X"00000020000000200000002000000020", 
10045=>X"00000020000000200000002000000020", 10046=>X"00000020000000200000002000000020", 10047=>X"00000020000000200000002000000020", 10048=>X"00000020000000200000002000000020", 10049=>X"00000020000000200000002000000020", 
10050=>X"00000020000000200000002000000020", 10051=>X"00000020000000200000002000000020", 10052=>X"00000020000000200000002000000020", 10053=>X"00000020000000200000002000000020", 10054=>X"00000020000000200000002000000020", 
10055=>X"00000020000000200000002000000020", 10056=>X"00000020000000200000002000000020", 10057=>X"00000020000000200000002000000020", 10058=>X"00000020000000200000002000000020", 10059=>X"00000020000000200000002000000020", 
10060=>X"00000020000000200000002000000020", 10061=>X"00000020000000200000002000000020", 10062=>X"00000020000000200000002000000020", 10063=>X"00000020000000200000002000000020", 10064=>X"00000020000000200000002000000020", 
10065=>X"00000020000000200000002000000020", 10066=>X"00000020000000200000002000000020", 10067=>X"00000020000000200000002000000020", 10068=>X"00000020000000200000002000000020", 10069=>X"00000020000000200000002000000020", 
10070=>X"00000020000000200000002000000020", 10071=>X"00000020000000200000002000000020", 10072=>X"00000020000000200000002000000020", 10073=>X"00000020000000200000002000000020", 10074=>X"00000020000000200000002000000020", 
10075=>X"00000020000000200000002000000020", 10076=>X"00000020000000200000002000000020", 10077=>X"00000020000000200000002000000020", 10078=>X"00000020000000200000002000000020", 10079=>X"00000020000000200000002000000020", 
10080=>X"00000020000000200000002000000020", 10081=>X"00000020000000200000002000000020", 10082=>X"00000020000000200000002000000020", 10083=>X"00000020000000200000002000000020", 10084=>X"00000020000000200000002000000020", 
10085=>X"00000020000000200000002000000020", 10086=>X"00000020000000200000002000000020", 10087=>X"00000020000000200000002000000020", 10088=>X"00000020000000200000002000000020", 10089=>X"00000020000000200000002000000020", 
10090=>X"00000020000000200000002000000020", 10091=>X"00000020000000200000002000000020", 10092=>X"00000020000000200000002000000020", 10093=>X"00000020000000200000002000000020", 10094=>X"00000020000000200000002000000020", 
10095=>X"00000020000000200000002000000020", 10096=>X"00000020000000200000002000000020", 10097=>X"00000020000000200000002000000020", 10098=>X"00000020000000200000002000000020", 10099=>X"00000020000000200000002000000020", 
10100=>X"00000020000000200000002000000020", 10101=>X"00000020000000200000002000000020", 10102=>X"00000020000000200000002000000020", 10103=>X"00000020000000200000002000000020", 10104=>X"00000020000000200000002000000020", 
10105=>X"00000020000000200000002000000020", 10106=>X"00000020000000200000002000000020", 10107=>X"00000020000000200000002000000020", 10108=>X"00000020000000200000002000000020", 10109=>X"00000020000000200000002000000020", 
10110=>X"00000020000000200000002000000020", 10111=>X"00000020000000200000002000000020", 10112=>X"00000020000000200000002000000020", 10113=>X"00000020000000200000002000000020", 10114=>X"00000020000000200000002000000020", 
10115=>X"00000020000000200000002000000020", 10116=>X"00000020000000200000002000000020", 10117=>X"00000020000000200000002000000020", 10118=>X"00000020000000200000002000000020", 10119=>X"00000020000000200000002000000020", 
10120=>X"00000020000000200000002000000020", 10121=>X"00000020000000200000002000000020", 10122=>X"00000020000000200000002000000020", 10123=>X"00000020000000200000002000000020", 10124=>X"00000020000000200000002000000020", 
10125=>X"00000020000000200000002000000020", 10126=>X"00000020000000200000002000000020", 10127=>X"00000020000000200000002000000020", 10128=>X"00000020000000200000002000000020", 10129=>X"00000020000000200000002000000020", 
10130=>X"00000020000000200000002000000020", 10131=>X"00000020000000200000002000000020", 10132=>X"00000020000000200000002000000020", 10133=>X"00000020000000200000002000000020", 10134=>X"00000020000000200000002000000020", 
10135=>X"00000020000000200000002000000020", 10136=>X"00000020000000200000002000000020", 10137=>X"00000020000000200000002000000020", 10138=>X"00000020000000200000002000000020", 10139=>X"00000020000000200000002000000020", 
10140=>X"00000020000000200000002000000020", 10141=>X"00000020000000200000002000000020", 10142=>X"00000020000000200000002000000020", 10143=>X"00000020000000200000002000000020", 10144=>X"00000020000000200000002000000020", 
10145=>X"00000020000000200000002000000020", 10146=>X"00000020000000200000002000000020", 10147=>X"00000020000000200000002000000020", 10148=>X"00000020000000200000002000000020", 10149=>X"00000020000000200000002000000020", 
10150=>X"00000020000000200000002000000020", 10151=>X"00000020000000200000002000000020", 10152=>X"00000020000000200000002000000020", 10153=>X"00000020000000200000002000000020", 10154=>X"00000020000000200000002000000020", 
10155=>X"00000020000000200000002000000020", 10156=>X"00000020000000200000002000000020", 10157=>X"00000020000000200000002000000020", 10158=>X"00000020000000200000002000000020", 10159=>X"00000020000000200000002000000020", 
10160=>X"00000020000000200000002000000020", 10161=>X"00000020000000200000002000000020", 10162=>X"00000020000000200000002000000020", 10163=>X"00000020000000200000002000000020", 10164=>X"00000020000000200000002000000020", 
10165=>X"00000020000000200000002000000020", 10166=>X"00000020000000200000002000000020", 10167=>X"00000020000000200000002000000020", 10168=>X"00000020000000200000002000000020", 10169=>X"00000020000000200000002000000020", 
10170=>X"00000020000000200000002000000020", 10171=>X"00000020000000200000002000000020", 10172=>X"00000020000000200000002000000020", 10173=>X"00000020000000200000002000000020", 10174=>X"00000020000000200000002000000020", 
10175=>X"00000020000000200000002000000020", 10176=>X"00000020000000200000002000000020", 10177=>X"00000020000000200000002000000020", 10178=>X"00000020000000200000002000000020", 10179=>X"00000020000000200000002000000020", 
10180=>X"00000020000000200000002000000020", 10181=>X"00000020000000200000002000000020", 10182=>X"00000020000000200000002000000020", 10183=>X"00000020000000200000002000000020", 10184=>X"00000020000000200000002000000020", 
10185=>X"00000020000000200000002000000020", 10186=>X"00000020000000200000002000000020", 10187=>X"00000020000000200000002000000020", 10188=>X"00000020000000200000002000000020", 10189=>X"00000020000000200000002000000020", 
10190=>X"00000020000000200000002000000020", 10191=>X"00000020000000200000002000000020", 10192=>X"0000001f0000001f0000001f0000001f", 10193=>X"0000001f0000001f0000001f0000001f", 10194=>X"0000001f0000001f0000001f0000001f", 
10195=>X"0000001f0000001f0000001f0000001f", 10196=>X"0000001f0000001f0000001f0000001f", 10197=>X"0000001f0000001f0000001f0000001f", 10198=>X"0000001f0000001f0000001f0000001f", 10199=>X"0000001f0000001f0000001f0000001f", 
10200=>X"0000001f0000001f0000001f0000001f", 10201=>X"0000001f0000001f0000001f0000001f", 10202=>X"0000001f0000001f0000001f0000001f", 10203=>X"0000001f0000001f0000001f0000001f", 10204=>X"0000001f0000001f0000001f0000001f", 
10205=>X"0000001f0000001f0000001f0000001f", 10206=>X"0000001f0000001f0000001f0000001f", 10207=>X"0000001f0000001f0000001f0000001f", 10208=>X"0000001f0000001f0000001f0000001f", 10209=>X"0000001f0000001f0000001f0000001f", 
10210=>X"0000001f0000001f0000001f0000001f", 10211=>X"0000001f0000001f0000001f0000001f", 10212=>X"0000001f0000001f0000001f0000001f", 10213=>X"0000001f0000001f0000001f0000001f", 10214=>X"0000001f0000001f0000001f0000001f", 
10215=>X"0000001f0000001f0000001f0000001f", 10216=>X"0000001f0000001f0000001f0000001f", 10217=>X"0000001f0000001f0000001f0000001f", 10218=>X"0000001f0000001f0000001f0000001f", 10219=>X"0000001f0000001f0000001f0000001f", 
10220=>X"0000001f0000001f0000001f0000001f", 10221=>X"0000001f0000001f0000001f0000001f", 10222=>X"0000001f0000001f0000001f0000001f", 10223=>X"0000001f0000001f0000001f0000001f", 10224=>X"0000001f0000001f0000001f0000001f", 
10225=>X"0000001f0000001f0000001f0000001f", 10226=>X"0000001f0000001f0000001f0000001f", 10227=>X"0000001f0000001f0000001f0000001f", 10228=>X"0000001f0000001f0000001f0000001f", 10229=>X"0000001f0000001f0000001f0000001f", 
10230=>X"0000001f0000001f0000001f0000001f", 10231=>X"0000001f0000001f0000001f0000001f", 10232=>X"0000001f0000001f0000001f0000001f", 10233=>X"0000001f0000001f0000001f0000001f", 10234=>X"0000001f0000001f0000001f0000001f", 
10235=>X"0000001f0000001f0000001f0000001f", 10236=>X"0000001f0000001f0000001f0000001f", 10237=>X"0000001f0000001f0000001f0000001f", 10238=>X"0000001f0000001f0000001f0000001f", 10239=>X"0000001f0000001f0000001f0000001f", 
10240=>X"0000001f0000001f0000001f0000001f", 10241=>X"0000001f0000001f0000001f0000001f", 10242=>X"0000001f0000001f0000001f0000001f", 10243=>X"0000001f0000001f0000001f0000001f", 10244=>X"0000001f0000001f0000001f0000001f", 
10245=>X"0000001f0000001f0000001f0000001f", 10246=>X"0000001f0000001f0000001f0000001f", 10247=>X"0000001f0000001f0000001f0000001f", 10248=>X"0000001f0000001f0000001f0000001f", 10249=>X"0000001f0000001f0000001f0000001f", 
10250=>X"0000001f0000001f0000001f0000001f", 10251=>X"0000001f0000001f0000001f0000001f", 10252=>X"0000001f0000001f0000001f0000001f", 10253=>X"0000001f0000001f0000001f0000001f", 10254=>X"0000001f0000001f0000001f0000001f", 
10255=>X"0000001f0000001f0000001f0000001f", 10256=>X"0000001f0000001f0000001f0000001f", 10257=>X"0000001f0000001f0000001f0000001f", 10258=>X"0000001f0000001f0000001f0000001f", 10259=>X"0000001f0000001f0000001f0000001f", 
10260=>X"0000001f0000001f0000001f0000001f", 10261=>X"0000001f0000001f0000001f0000001f", 10262=>X"0000001f0000001f0000001f0000001f", 10263=>X"0000001f0000001f0000001f0000001f", 10264=>X"0000001f0000001f0000001f0000001f", 
10265=>X"0000001f0000001f0000001f0000001f", 10266=>X"0000001f0000001f0000001f0000001f", 10267=>X"0000001f0000001f0000001f0000001f", 10268=>X"0000001f0000001f0000001f0000001f", 10269=>X"0000001f0000001f0000001f0000001f", 
10270=>X"0000001f0000001f0000001f0000001f", 10271=>X"0000001f0000001f0000001f0000001f", 10272=>X"0000001f0000001f0000001f0000001f", 10273=>X"0000001f0000001f0000001f0000001f", 10274=>X"0000001f0000001f0000001f0000001f", 
10275=>X"0000001f0000001f0000001f0000001f", 10276=>X"0000001f0000001f0000001f0000001f", 10277=>X"0000001f0000001f0000001f0000001f", 10278=>X"0000001f0000001f0000001f0000001f", 10279=>X"0000001f0000001f0000001f0000001f", 
10280=>X"0000001f0000001f0000001f0000001f", 10281=>X"0000001f0000001f0000001f0000001f", 10282=>X"0000001f0000001f0000001f0000001f", 10283=>X"0000001f0000001f0000001f0000001f", 10284=>X"0000001f0000001f0000001f0000001f", 
10285=>X"0000001f0000001f0000001f0000001f", 10286=>X"0000001f0000001f0000001f0000001f", 10287=>X"0000001f0000001f0000001f0000001f", 10288=>X"0000001f0000001f0000001f0000001f", 10289=>X"0000001f0000001f0000001f0000001f", 
10290=>X"0000001f0000001f0000001f0000001f", 10291=>X"0000001f0000001f0000001f0000001f", 10292=>X"0000001f0000001f0000001f0000001f", 10293=>X"0000001f0000001f0000001f0000001f", 10294=>X"0000001f0000001f0000001f0000001f", 
10295=>X"0000001f0000001f0000001f0000001f", 10296=>X"0000001f0000001f0000001f0000001f", 10297=>X"0000001f0000001f0000001f0000001f", 10298=>X"0000001f0000001f0000001f0000001f", 10299=>X"0000001f0000001f0000001f0000001f", 
10300=>X"0000001f0000001f0000001f0000001f", 10301=>X"0000001f0000001f0000001f0000001f", 10302=>X"0000001f0000001f0000001f0000001f", 10303=>X"0000001f0000001f0000001f0000001f", 10304=>X"0000001f0000001f0000001f0000001f", 
10305=>X"0000001f0000001f0000001f0000001f", 10306=>X"0000001f0000001f0000001f0000001f", 10307=>X"0000001f0000001f0000001f0000001f", 10308=>X"0000001f0000001f0000001f0000001f", 10309=>X"0000001f0000001f0000001f0000001f", 
10310=>X"0000001f0000001f0000001f0000001f", 10311=>X"0000001f0000001f0000001f0000001f", 10312=>X"0000001f0000001f0000001f0000001f", 10313=>X"0000001f0000001f0000001f0000001f", 10314=>X"0000001f0000001f0000001f0000001f", 
10315=>X"0000001f0000001f0000001f0000001f", 10316=>X"0000001f0000001f0000001f0000001f", 10317=>X"0000001f0000001f0000001f0000001f", 10318=>X"0000001f0000001f0000001f0000001f", 10319=>X"0000001f0000001f0000001f0000001f", 
10320=>X"0000001f0000001f0000001f0000001f", 10321=>X"0000001f0000001f0000001f0000001f", 10322=>X"0000001f0000001f0000001f0000001f", 10323=>X"0000001f0000001f0000001f0000001f", 10324=>X"0000001f0000001f0000001f0000001f", 
10325=>X"0000001f0000001f0000001f0000001f", 10326=>X"0000001f0000001f0000001f0000001f", 10327=>X"0000001f0000001f0000001f0000001f", 10328=>X"0000001f0000001f0000001f0000001f", 10329=>X"0000001f0000001f0000001f0000001f", 
10330=>X"0000001f0000001f0000001f0000001f", 10331=>X"0000001f0000001f0000001f0000001f", 10332=>X"0000001f0000001f0000001f0000001f", 10333=>X"0000001f0000001f0000001f0000001f", 10334=>X"0000001f0000001f0000001f0000001f", 
10335=>X"0000001f0000001f0000001f0000001f", 10336=>X"0000001f0000001f0000001f0000001f", 10337=>X"0000001f0000001f0000001f0000001f", 10338=>X"0000001f0000001f0000001f0000001f", 10339=>X"0000001f0000001f0000001f0000001f", 
10340=>X"0000001f0000001f0000001f0000001f", 10341=>X"0000001f0000001f0000001f0000001f", 10342=>X"0000001f0000001f0000001f0000001f", 10343=>X"0000001f0000001f0000001f0000001f", 10344=>X"0000001f0000001f0000001f0000001f", 
10345=>X"0000001f0000001f0000001f0000001f", 10346=>X"0000001f0000001f0000001f0000001f", 10347=>X"0000001f0000001f0000001f0000001f", 10348=>X"0000001f0000001f0000001f0000001f", 10349=>X"0000001f0000001f0000001f0000001f", 
10350=>X"0000001f0000001f0000001f0000001f", 10351=>X"0000001f0000001f0000001f0000001f", 10352=>X"0000001f0000001f0000001f0000001f", 10353=>X"0000001f0000001f0000001f0000001f", 10354=>X"0000001f0000001f0000001f0000001f", 
10355=>X"0000001f0000001f0000001f0000001f", 10356=>X"0000001f0000001f0000001f0000001f", 10357=>X"0000001f0000001f0000001f0000001f", 10358=>X"0000001f0000001f0000001f0000001f", 10359=>X"0000001f0000001f0000001f0000001f", 
10360=>X"0000001f0000001f0000001f0000001f", 10361=>X"0000001f0000001f0000001f0000001f", 10362=>X"0000001f0000001f0000001f0000001f", 10363=>X"0000001f0000001f0000001f0000001f", 10364=>X"0000001f0000001f0000001f0000001f", 
10365=>X"0000001f0000001f0000001f0000001f", 10366=>X"0000001f0000001f0000001f0000001f", 10367=>X"0000001f0000001f0000001f0000001f", 10368=>X"0000001f0000001f0000001f0000001f", 10369=>X"0000001f0000001f0000001f0000001f", 
10370=>X"0000001f0000001f0000001f0000001f", 10371=>X"0000001f0000001f0000001f0000001f", 10372=>X"0000001f0000001f0000001f0000001f", 10373=>X"0000001f0000001f0000001f0000001f", 10374=>X"0000001f0000001f0000001f0000001f", 
10375=>X"0000001f0000001f0000001f0000001f", 10376=>X"0000001f0000001f0000001f0000001f", 10377=>X"0000001f0000001f0000001f0000001f", 10378=>X"0000001f0000001f0000001f0000001f", 10379=>X"0000001f0000001f0000001f0000001f", 
10380=>X"0000001f0000001f0000001f0000001f", 10381=>X"0000001f0000001f0000001f0000001f", 10382=>X"0000001f0000001f0000001f0000001f", 10383=>X"0000001f0000001f0000001f0000001f", 10384=>X"0000001f0000001f0000001f0000001f", 
10385=>X"0000001f0000001f0000001f0000001f", 10386=>X"0000001f0000001f0000001f0000001f", 10387=>X"0000001f0000001f0000001f0000001f", 10388=>X"0000001f0000001f0000001f0000001f", 10389=>X"0000001f0000001f0000001f0000001f", 
10390=>X"0000001f0000001f0000001f0000001f", 10391=>X"0000001f0000001f0000001f0000001f", 10392=>X"0000001f0000001f0000001f0000001f", 10393=>X"0000001f0000001f0000001f0000001f", 10394=>X"0000001f0000001f0000001f0000001f", 
10395=>X"0000001f0000001f0000001f0000001f", 10396=>X"0000001f0000001f0000001f0000001f", 10397=>X"0000001f0000001f0000001f0000001f", 10398=>X"0000001f0000001f0000001f0000001f", 10399=>X"0000001f0000001f0000001f0000001f", 
10400=>X"0000001f0000001f0000001f0000001f", 10401=>X"0000001f0000001f0000001f0000001f", 10402=>X"0000001f0000001f0000001f0000001f", 10403=>X"0000001f0000001f0000001f0000001f", 10404=>X"0000001f0000001f0000001f0000001f", 
10405=>X"0000001f0000001f0000001f0000001f", 10406=>X"0000001f0000001f0000001f0000001f", 10407=>X"0000001f0000001f0000001f0000001f", 10408=>X"0000001f0000001f0000001f0000001f", 10409=>X"0000001f0000001f0000001f0000001f", 
10410=>X"0000001f0000001f0000001f0000001f", 10411=>X"0000001f0000001f0000001f0000001f", 10412=>X"0000001f0000001f0000001f0000001f", 10413=>X"0000001f0000001f0000001f0000001f", 10414=>X"0000001f0000001f0000001f0000001f", 
10415=>X"0000001f0000001f0000001f0000001f", 10416=>X"0000001f0000001f0000001f0000001f", 10417=>X"0000001f0000001f0000001f0000001f", 10418=>X"0000001f0000001f0000001f0000001f", 10419=>X"0000001f0000001f0000001f0000001f", 
10420=>X"0000001f0000001f0000001f0000001f", 10421=>X"0000001f0000001f0000001f0000001f", 10422=>X"0000001f0000001f0000001f0000001f", 10423=>X"0000001f0000001f0000001f0000001f", 10424=>X"0000001f0000001f0000001f0000001f", 
10425=>X"0000001f0000001f0000001f0000001f", 10426=>X"0000001f0000001f0000001f0000001f", 10427=>X"0000001f0000001f0000001f0000001f", 10428=>X"0000001f0000001f0000001f0000001f", 10429=>X"0000001f0000001f0000001f0000001f", 
10430=>X"0000001f0000001f0000001f0000001f", 10431=>X"0000001f0000001f0000001f0000001f", 10432=>X"0000001f0000001f0000001f0000001f", 10433=>X"0000001f0000001f0000001f0000001f", 10434=>X"0000001f0000001f0000001f0000001f", 
10435=>X"0000001f0000001f0000001f0000001f", 10436=>X"0000001f0000001f0000001f0000001f", 10437=>X"0000001f0000001f0000001f0000001f", 10438=>X"0000001f0000001f0000001f0000001f", 10439=>X"0000001f0000001f0000001f0000001f", 
10440=>X"0000001f0000001f0000001f0000001f", 10441=>X"0000001f0000001f0000001f0000001f", 10442=>X"0000001f0000001f0000001f0000001f", 10443=>X"0000001f0000001f0000001f0000001f", 10444=>X"0000001f0000001f0000001f0000001f", 
10445=>X"0000001f0000001f0000001f0000001f", 10446=>X"0000001f0000001f0000001f0000001f", 10447=>X"0000001f0000001f0000001f0000001f", 10448=>X"0000001f0000001f0000001f0000001f", 10449=>X"0000001f0000001f0000001f0000001f", 
10450=>X"0000001f0000001f0000001f0000001f", 10451=>X"0000001f0000001f0000001f0000001f", 10452=>X"0000001f0000001f0000001f0000001f", 10453=>X"0000001f0000001f0000001f0000001f", 10454=>X"0000001f0000001f0000001f0000001f", 
10455=>X"0000001f0000001f0000001f0000001f", 10456=>X"0000001f0000001f0000001f0000001f", 10457=>X"0000001f0000001f0000001f0000001f", 10458=>X"0000001f0000001f0000001f0000001f", 10459=>X"0000001f0000001f0000001f0000001f", 
10460=>X"0000001f0000001f0000001f0000001f", 10461=>X"0000001f0000001f0000001f0000001f", 10462=>X"0000001f0000001f0000001f0000001f", 10463=>X"0000001f0000001f0000001f0000001f", 10464=>X"0000001e0000001f0000001f0000001f", 
10465=>X"0000001e0000001e0000001e0000001e", 10466=>X"0000001e0000001e0000001e0000001e", 10467=>X"0000001e0000001e0000001e0000001e", 10468=>X"0000001e0000001e0000001e0000001e", 10469=>X"0000001e0000001e0000001e0000001e", 
10470=>X"0000001e0000001e0000001e0000001e", 10471=>X"0000001e0000001e0000001e0000001e", 10472=>X"0000001e0000001e0000001e0000001e", 10473=>X"0000001e0000001e0000001e0000001e", 10474=>X"0000001e0000001e0000001e0000001e", 
10475=>X"0000001e0000001e0000001e0000001e", 10476=>X"0000001e0000001e0000001e0000001e", 10477=>X"0000001e0000001e0000001e0000001e", 10478=>X"0000001e0000001e0000001e0000001e", 10479=>X"0000001e0000001e0000001e0000001e", 
10480=>X"0000001e0000001e0000001e0000001e", 10481=>X"0000001e0000001e0000001e0000001e", 10482=>X"0000001e0000001e0000001e0000001e", 10483=>X"0000001e0000001e0000001e0000001e", 10484=>X"0000001e0000001e0000001e0000001e", 
10485=>X"0000001e0000001e0000001e0000001e", 10486=>X"0000001e0000001e0000001e0000001e", 10487=>X"0000001e0000001e0000001e0000001e", 10488=>X"0000001e0000001e0000001e0000001e", 10489=>X"0000001e0000001e0000001e0000001e", 
10490=>X"0000001e0000001e0000001e0000001e", 10491=>X"0000001e0000001e0000001e0000001e", 10492=>X"0000001e0000001e0000001e0000001e", 10493=>X"0000001e0000001e0000001e0000001e", 10494=>X"0000001e0000001e0000001e0000001e", 
10495=>X"0000001e0000001e0000001e0000001e", 10496=>X"0000001e0000001e0000001e0000001e", 10497=>X"0000001e0000001e0000001e0000001e", 10498=>X"0000001e0000001e0000001e0000001e", 10499=>X"0000001e0000001e0000001e0000001e", 
10500=>X"0000001e0000001e0000001e0000001e", 10501=>X"0000001e0000001e0000001e0000001e", 10502=>X"0000001e0000001e0000001e0000001e", 10503=>X"0000001e0000001e0000001e0000001e", 10504=>X"0000001e0000001e0000001e0000001e", 
10505=>X"0000001e0000001e0000001e0000001e", 10506=>X"0000001e0000001e0000001e0000001e", 10507=>X"0000001e0000001e0000001e0000001e", 10508=>X"0000001e0000001e0000001e0000001e", 10509=>X"0000001e0000001e0000001e0000001e", 
10510=>X"0000001e0000001e0000001e0000001e", 10511=>X"0000001e0000001e0000001e0000001e", 10512=>X"0000001e0000001e0000001e0000001e", 10513=>X"0000001e0000001e0000001e0000001e", 10514=>X"0000001e0000001e0000001e0000001e", 
10515=>X"0000001e0000001e0000001e0000001e", 10516=>X"0000001e0000001e0000001e0000001e", 10517=>X"0000001e0000001e0000001e0000001e", 10518=>X"0000001e0000001e0000001e0000001e", 10519=>X"0000001e0000001e0000001e0000001e", 
10520=>X"0000001e0000001e0000001e0000001e", 10521=>X"0000001e0000001e0000001e0000001e", 10522=>X"0000001e0000001e0000001e0000001e", 10523=>X"0000001e0000001e0000001e0000001e", 10524=>X"0000001e0000001e0000001e0000001e", 
10525=>X"0000001e0000001e0000001e0000001e", 10526=>X"0000001e0000001e0000001e0000001e", 10527=>X"0000001e0000001e0000001e0000001e", 10528=>X"0000001e0000001e0000001e0000001e", 10529=>X"0000001e0000001e0000001e0000001e", 
10530=>X"0000001e0000001e0000001e0000001e", 10531=>X"0000001e0000001e0000001e0000001e", 10532=>X"0000001e0000001e0000001e0000001e", 10533=>X"0000001e0000001e0000001e0000001e", 10534=>X"0000001e0000001e0000001e0000001e", 
10535=>X"0000001e0000001e0000001e0000001e", 10536=>X"0000001e0000001e0000001e0000001e", 10537=>X"0000001e0000001e0000001e0000001e", 10538=>X"0000001e0000001e0000001e0000001e", 10539=>X"0000001e0000001e0000001e0000001e", 
10540=>X"0000001e0000001e0000001e0000001e", 10541=>X"0000001e0000001e0000001e0000001e", 10542=>X"0000001e0000001e0000001e0000001e", 10543=>X"0000001e0000001e0000001e0000001e", 10544=>X"0000001e0000001e0000001e0000001e", 
10545=>X"0000001e0000001e0000001e0000001e", 10546=>X"0000001e0000001e0000001e0000001e", 10547=>X"0000001e0000001e0000001e0000001e", 10548=>X"0000001e0000001e0000001e0000001e", 10549=>X"0000001e0000001e0000001e0000001e", 
10550=>X"0000001e0000001e0000001e0000001e", 10551=>X"0000001e0000001e0000001e0000001e", 10552=>X"0000001e0000001e0000001e0000001e", 10553=>X"0000001e0000001e0000001e0000001e", 10554=>X"0000001e0000001e0000001e0000001e", 
10555=>X"0000001e0000001e0000001e0000001e", 10556=>X"0000001e0000001e0000001e0000001e", 10557=>X"0000001e0000001e0000001e0000001e", 10558=>X"0000001e0000001e0000001e0000001e", 10559=>X"0000001e0000001e0000001e0000001e", 
10560=>X"0000001e0000001e0000001e0000001e", 10561=>X"0000001e0000001e0000001e0000001e", 10562=>X"0000001e0000001e0000001e0000001e", 10563=>X"0000001e0000001e0000001e0000001e", 10564=>X"0000001e0000001e0000001e0000001e", 
10565=>X"0000001e0000001e0000001e0000001e", 10566=>X"0000001e0000001e0000001e0000001e", 10567=>X"0000001e0000001e0000001e0000001e", 10568=>X"0000001e0000001e0000001e0000001e", 10569=>X"0000001e0000001e0000001e0000001e", 
10570=>X"0000001e0000001e0000001e0000001e", 10571=>X"0000001e0000001e0000001e0000001e", 10572=>X"0000001e0000001e0000001e0000001e", 10573=>X"0000001e0000001e0000001e0000001e", 10574=>X"0000001e0000001e0000001e0000001e", 
10575=>X"0000001e0000001e0000001e0000001e", 10576=>X"0000001e0000001e0000001e0000001e", 10577=>X"0000001e0000001e0000001e0000001e", 10578=>X"0000001e0000001e0000001e0000001e", 10579=>X"0000001e0000001e0000001e0000001e", 
10580=>X"0000001e0000001e0000001e0000001e", 10581=>X"0000001e0000001e0000001e0000001e", 10582=>X"0000001e0000001e0000001e0000001e", 10583=>X"0000001e0000001e0000001e0000001e", 10584=>X"0000001e0000001e0000001e0000001e", 
10585=>X"0000001e0000001e0000001e0000001e", 10586=>X"0000001e0000001e0000001e0000001e", 10587=>X"0000001e0000001e0000001e0000001e", 10588=>X"0000001e0000001e0000001e0000001e", 10589=>X"0000001e0000001e0000001e0000001e", 
10590=>X"0000001e0000001e0000001e0000001e", 10591=>X"0000001e0000001e0000001e0000001e", 10592=>X"0000001e0000001e0000001e0000001e", 10593=>X"0000001e0000001e0000001e0000001e", 10594=>X"0000001e0000001e0000001e0000001e", 
10595=>X"0000001e0000001e0000001e0000001e", 10596=>X"0000001e0000001e0000001e0000001e", 10597=>X"0000001e0000001e0000001e0000001e", 10598=>X"0000001e0000001e0000001e0000001e", 10599=>X"0000001e0000001e0000001e0000001e", 
10600=>X"0000001e0000001e0000001e0000001e", 10601=>X"0000001e0000001e0000001e0000001e", 10602=>X"0000001e0000001e0000001e0000001e", 10603=>X"0000001e0000001e0000001e0000001e", 10604=>X"0000001e0000001e0000001e0000001e", 
10605=>X"0000001e0000001e0000001e0000001e", 10606=>X"0000001e0000001e0000001e0000001e", 10607=>X"0000001e0000001e0000001e0000001e", 10608=>X"0000001e0000001e0000001e0000001e", 10609=>X"0000001e0000001e0000001e0000001e", 
10610=>X"0000001e0000001e0000001e0000001e", 10611=>X"0000001e0000001e0000001e0000001e", 10612=>X"0000001e0000001e0000001e0000001e", 10613=>X"0000001e0000001e0000001e0000001e", 10614=>X"0000001e0000001e0000001e0000001e", 
10615=>X"0000001e0000001e0000001e0000001e", 10616=>X"0000001e0000001e0000001e0000001e", 10617=>X"0000001e0000001e0000001e0000001e", 10618=>X"0000001e0000001e0000001e0000001e", 10619=>X"0000001e0000001e0000001e0000001e", 
10620=>X"0000001e0000001e0000001e0000001e", 10621=>X"0000001e0000001e0000001e0000001e", 10622=>X"0000001e0000001e0000001e0000001e", 10623=>X"0000001e0000001e0000001e0000001e", 10624=>X"0000001e0000001e0000001e0000001e", 
10625=>X"0000001e0000001e0000001e0000001e", 10626=>X"0000001e0000001e0000001e0000001e", 10627=>X"0000001e0000001e0000001e0000001e", 10628=>X"0000001e0000001e0000001e0000001e", 10629=>X"0000001e0000001e0000001e0000001e", 
10630=>X"0000001e0000001e0000001e0000001e", 10631=>X"0000001e0000001e0000001e0000001e", 10632=>X"0000001e0000001e0000001e0000001e", 10633=>X"0000001e0000001e0000001e0000001e", 10634=>X"0000001e0000001e0000001e0000001e", 
10635=>X"0000001e0000001e0000001e0000001e", 10636=>X"0000001e0000001e0000001e0000001e", 10637=>X"0000001e0000001e0000001e0000001e", 10638=>X"0000001e0000001e0000001e0000001e", 10639=>X"0000001e0000001e0000001e0000001e", 
10640=>X"0000001e0000001e0000001e0000001e", 10641=>X"0000001e0000001e0000001e0000001e", 10642=>X"0000001e0000001e0000001e0000001e", 10643=>X"0000001e0000001e0000001e0000001e", 10644=>X"0000001e0000001e0000001e0000001e", 
10645=>X"0000001e0000001e0000001e0000001e", 10646=>X"0000001e0000001e0000001e0000001e", 10647=>X"0000001e0000001e0000001e0000001e", 10648=>X"0000001e0000001e0000001e0000001e", 10649=>X"0000001e0000001e0000001e0000001e", 
10650=>X"0000001e0000001e0000001e0000001e", 10651=>X"0000001e0000001e0000001e0000001e", 10652=>X"0000001e0000001e0000001e0000001e", 10653=>X"0000001e0000001e0000001e0000001e", 10654=>X"0000001e0000001e0000001e0000001e", 
10655=>X"0000001e0000001e0000001e0000001e", 10656=>X"0000001e0000001e0000001e0000001e", 10657=>X"0000001e0000001e0000001e0000001e", 10658=>X"0000001e0000001e0000001e0000001e", 10659=>X"0000001e0000001e0000001e0000001e", 
10660=>X"0000001e0000001e0000001e0000001e", 10661=>X"0000001e0000001e0000001e0000001e", 10662=>X"0000001e0000001e0000001e0000001e", 10663=>X"0000001e0000001e0000001e0000001e", 10664=>X"0000001e0000001e0000001e0000001e", 
10665=>X"0000001e0000001e0000001e0000001e", 10666=>X"0000001e0000001e0000001e0000001e", 10667=>X"0000001e0000001e0000001e0000001e", 10668=>X"0000001e0000001e0000001e0000001e", 10669=>X"0000001e0000001e0000001e0000001e", 
10670=>X"0000001e0000001e0000001e0000001e", 10671=>X"0000001e0000001e0000001e0000001e", 10672=>X"0000001e0000001e0000001e0000001e", 10673=>X"0000001e0000001e0000001e0000001e", 10674=>X"0000001e0000001e0000001e0000001e", 
10675=>X"0000001e0000001e0000001e0000001e", 10676=>X"0000001e0000001e0000001e0000001e", 10677=>X"0000001e0000001e0000001e0000001e", 10678=>X"0000001e0000001e0000001e0000001e", 10679=>X"0000001e0000001e0000001e0000001e", 
10680=>X"0000001e0000001e0000001e0000001e", 10681=>X"0000001e0000001e0000001e0000001e", 10682=>X"0000001e0000001e0000001e0000001e", 10683=>X"0000001e0000001e0000001e0000001e", 10684=>X"0000001e0000001e0000001e0000001e", 
10685=>X"0000001e0000001e0000001e0000001e", 10686=>X"0000001e0000001e0000001e0000001e", 10687=>X"0000001e0000001e0000001e0000001e", 10688=>X"0000001e0000001e0000001e0000001e", 10689=>X"0000001e0000001e0000001e0000001e", 
10690=>X"0000001e0000001e0000001e0000001e", 10691=>X"0000001e0000001e0000001e0000001e", 10692=>X"0000001e0000001e0000001e0000001e", 10693=>X"0000001e0000001e0000001e0000001e", 10694=>X"0000001e0000001e0000001e0000001e", 
10695=>X"0000001e0000001e0000001e0000001e", 10696=>X"0000001e0000001e0000001e0000001e", 10697=>X"0000001e0000001e0000001e0000001e", 10698=>X"0000001e0000001e0000001e0000001e", 10699=>X"0000001e0000001e0000001e0000001e", 
10700=>X"0000001e0000001e0000001e0000001e", 10701=>X"0000001e0000001e0000001e0000001e", 10702=>X"0000001e0000001e0000001e0000001e", 10703=>X"0000001e0000001e0000001e0000001e", 10704=>X"0000001e0000001e0000001e0000001e", 
10705=>X"0000001e0000001e0000001e0000001e", 10706=>X"0000001e0000001e0000001e0000001e", 10707=>X"0000001e0000001e0000001e0000001e", 10708=>X"0000001e0000001e0000001e0000001e", 10709=>X"0000001e0000001e0000001e0000001e", 
10710=>X"0000001e0000001e0000001e0000001e", 10711=>X"0000001e0000001e0000001e0000001e", 10712=>X"0000001e0000001e0000001e0000001e", 10713=>X"0000001e0000001e0000001e0000001e", 10714=>X"0000001e0000001e0000001e0000001e", 
10715=>X"0000001e0000001e0000001e0000001e", 10716=>X"0000001e0000001e0000001e0000001e", 10717=>X"0000001e0000001e0000001e0000001e", 10718=>X"0000001e0000001e0000001e0000001e", 10719=>X"0000001e0000001e0000001e0000001e", 
10720=>X"0000001e0000001e0000001e0000001e", 10721=>X"0000001e0000001e0000001e0000001e", 10722=>X"0000001e0000001e0000001e0000001e", 10723=>X"0000001e0000001e0000001e0000001e", 10724=>X"0000001e0000001e0000001e0000001e", 
10725=>X"0000001e0000001e0000001e0000001e", 10726=>X"0000001e0000001e0000001e0000001e", 10727=>X"0000001e0000001e0000001e0000001e", 10728=>X"0000001e0000001e0000001e0000001e", 10729=>X"0000001e0000001e0000001e0000001e", 
10730=>X"0000001e0000001e0000001e0000001e", 10731=>X"0000001e0000001e0000001e0000001e", 10732=>X"0000001e0000001e0000001e0000001e", 10733=>X"0000001e0000001e0000001e0000001e", 10734=>X"0000001e0000001e0000001e0000001e", 
10735=>X"0000001e0000001e0000001e0000001e", 10736=>X"0000001e0000001e0000001e0000001e", 10737=>X"0000001e0000001e0000001e0000001e", 10738=>X"0000001e0000001e0000001e0000001e", 10739=>X"0000001e0000001e0000001e0000001e", 
10740=>X"0000001e0000001e0000001e0000001e", 10741=>X"0000001e0000001e0000001e0000001e", 10742=>X"0000001e0000001e0000001e0000001e", 10743=>X"0000001e0000001e0000001e0000001e", 10744=>X"0000001e0000001e0000001e0000001e", 
10745=>X"0000001e0000001e0000001e0000001e", 10746=>X"0000001e0000001e0000001e0000001e", 10747=>X"0000001e0000001e0000001e0000001e", 10748=>X"0000001e0000001e0000001e0000001e", 10749=>X"0000001e0000001e0000001e0000001e", 
10750=>X"0000001e0000001e0000001e0000001e", 10751=>X"0000001e0000001e0000001e0000001e", 10752=>X"0000001e0000001e0000001e0000001e", 10753=>X"0000001e0000001e0000001e0000001e", 10754=>X"0000001e0000001e0000001e0000001e", 
10755=>X"0000001e0000001e0000001e0000001e", 10756=>X"0000001d0000001d0000001d0000001d", 10757=>X"0000001d0000001d0000001d0000001d", 10758=>X"0000001d0000001d0000001d0000001d", 10759=>X"0000001d0000001d0000001d0000001d", 
10760=>X"0000001d0000001d0000001d0000001d", 10761=>X"0000001d0000001d0000001d0000001d", 10762=>X"0000001d0000001d0000001d0000001d", 10763=>X"0000001d0000001d0000001d0000001d", 10764=>X"0000001d0000001d0000001d0000001d", 
10765=>X"0000001d0000001d0000001d0000001d", 10766=>X"0000001d0000001d0000001d0000001d", 10767=>X"0000001d0000001d0000001d0000001d", 10768=>X"0000001d0000001d0000001d0000001d", 10769=>X"0000001d0000001d0000001d0000001d", 
10770=>X"0000001d0000001d0000001d0000001d", 10771=>X"0000001d0000001d0000001d0000001d", 10772=>X"0000001d0000001d0000001d0000001d", 10773=>X"0000001d0000001d0000001d0000001d", 10774=>X"0000001d0000001d0000001d0000001d", 
10775=>X"0000001d0000001d0000001d0000001d", 10776=>X"0000001d0000001d0000001d0000001d", 10777=>X"0000001d0000001d0000001d0000001d", 10778=>X"0000001d0000001d0000001d0000001d", 10779=>X"0000001d0000001d0000001d0000001d", 
10780=>X"0000001d0000001d0000001d0000001d", 10781=>X"0000001d0000001d0000001d0000001d", 10782=>X"0000001d0000001d0000001d0000001d", 10783=>X"0000001d0000001d0000001d0000001d", 10784=>X"0000001d0000001d0000001d0000001d", 
10785=>X"0000001d0000001d0000001d0000001d", 10786=>X"0000001d0000001d0000001d0000001d", 10787=>X"0000001d0000001d0000001d0000001d", 10788=>X"0000001d0000001d0000001d0000001d", 10789=>X"0000001d0000001d0000001d0000001d", 
10790=>X"0000001d0000001d0000001d0000001d", 10791=>X"0000001d0000001d0000001d0000001d", 10792=>X"0000001d0000001d0000001d0000001d", 10793=>X"0000001d0000001d0000001d0000001d", 10794=>X"0000001d0000001d0000001d0000001d", 
10795=>X"0000001d0000001d0000001d0000001d", 10796=>X"0000001d0000001d0000001d0000001d", 10797=>X"0000001d0000001d0000001d0000001d", 10798=>X"0000001d0000001d0000001d0000001d", 10799=>X"0000001d0000001d0000001d0000001d", 
10800=>X"0000001d0000001d0000001d0000001d", 10801=>X"0000001d0000001d0000001d0000001d", 10802=>X"0000001d0000001d0000001d0000001d", 10803=>X"0000001d0000001d0000001d0000001d", 10804=>X"0000001d0000001d0000001d0000001d", 
10805=>X"0000001d0000001d0000001d0000001d", 10806=>X"0000001d0000001d0000001d0000001d", 10807=>X"0000001d0000001d0000001d0000001d", 10808=>X"0000001d0000001d0000001d0000001d", 10809=>X"0000001d0000001d0000001d0000001d", 
10810=>X"0000001d0000001d0000001d0000001d", 10811=>X"0000001d0000001d0000001d0000001d", 10812=>X"0000001d0000001d0000001d0000001d", 10813=>X"0000001d0000001d0000001d0000001d", 10814=>X"0000001d0000001d0000001d0000001d", 
10815=>X"0000001d0000001d0000001d0000001d", 10816=>X"0000001d0000001d0000001d0000001d", 10817=>X"0000001d0000001d0000001d0000001d", 10818=>X"0000001d0000001d0000001d0000001d", 10819=>X"0000001d0000001d0000001d0000001d", 
10820=>X"0000001d0000001d0000001d0000001d", 10821=>X"0000001d0000001d0000001d0000001d", 10822=>X"0000001d0000001d0000001d0000001d", 10823=>X"0000001d0000001d0000001d0000001d", 10824=>X"0000001d0000001d0000001d0000001d", 
10825=>X"0000001d0000001d0000001d0000001d", 10826=>X"0000001d0000001d0000001d0000001d", 10827=>X"0000001d0000001d0000001d0000001d", 10828=>X"0000001d0000001d0000001d0000001d", 10829=>X"0000001d0000001d0000001d0000001d", 
10830=>X"0000001d0000001d0000001d0000001d", 10831=>X"0000001d0000001d0000001d0000001d", 10832=>X"0000001d0000001d0000001d0000001d", 10833=>X"0000001d0000001d0000001d0000001d", 10834=>X"0000001d0000001d0000001d0000001d", 
10835=>X"0000001d0000001d0000001d0000001d", 10836=>X"0000001d0000001d0000001d0000001d", 10837=>X"0000001d0000001d0000001d0000001d", 10838=>X"0000001d0000001d0000001d0000001d", 10839=>X"0000001d0000001d0000001d0000001d", 
10840=>X"0000001d0000001d0000001d0000001d", 10841=>X"0000001d0000001d0000001d0000001d", 10842=>X"0000001d0000001d0000001d0000001d", 10843=>X"0000001d0000001d0000001d0000001d", 10844=>X"0000001d0000001d0000001d0000001d", 
10845=>X"0000001d0000001d0000001d0000001d", 10846=>X"0000001d0000001d0000001d0000001d", 10847=>X"0000001d0000001d0000001d0000001d", 10848=>X"0000001d0000001d0000001d0000001d", 10849=>X"0000001d0000001d0000001d0000001d", 
10850=>X"0000001d0000001d0000001d0000001d", 10851=>X"0000001d0000001d0000001d0000001d", 10852=>X"0000001d0000001d0000001d0000001d", 10853=>X"0000001d0000001d0000001d0000001d", 10854=>X"0000001d0000001d0000001d0000001d", 
10855=>X"0000001d0000001d0000001d0000001d", 10856=>X"0000001d0000001d0000001d0000001d", 10857=>X"0000001d0000001d0000001d0000001d", 10858=>X"0000001d0000001d0000001d0000001d", 10859=>X"0000001d0000001d0000001d0000001d", 
10860=>X"0000001d0000001d0000001d0000001d", 10861=>X"0000001d0000001d0000001d0000001d", 10862=>X"0000001d0000001d0000001d0000001d", 10863=>X"0000001d0000001d0000001d0000001d", 10864=>X"0000001d0000001d0000001d0000001d", 
10865=>X"0000001d0000001d0000001d0000001d", 10866=>X"0000001d0000001d0000001d0000001d", 10867=>X"0000001d0000001d0000001d0000001d", 10868=>X"0000001d0000001d0000001d0000001d", 10869=>X"0000001d0000001d0000001d0000001d", 
10870=>X"0000001d0000001d0000001d0000001d", 10871=>X"0000001d0000001d0000001d0000001d", 10872=>X"0000001d0000001d0000001d0000001d", 10873=>X"0000001d0000001d0000001d0000001d", 10874=>X"0000001d0000001d0000001d0000001d", 
10875=>X"0000001d0000001d0000001d0000001d", 10876=>X"0000001d0000001d0000001d0000001d", 10877=>X"0000001d0000001d0000001d0000001d", 10878=>X"0000001d0000001d0000001d0000001d", 10879=>X"0000001d0000001d0000001d0000001d", 
10880=>X"0000001d0000001d0000001d0000001d", 10881=>X"0000001d0000001d0000001d0000001d", 10882=>X"0000001d0000001d0000001d0000001d", 10883=>X"0000001d0000001d0000001d0000001d", 10884=>X"0000001d0000001d0000001d0000001d", 
10885=>X"0000001d0000001d0000001d0000001d", 10886=>X"0000001d0000001d0000001d0000001d", 10887=>X"0000001d0000001d0000001d0000001d", 10888=>X"0000001d0000001d0000001d0000001d", 10889=>X"0000001d0000001d0000001d0000001d", 
10890=>X"0000001d0000001d0000001d0000001d", 10891=>X"0000001d0000001d0000001d0000001d", 10892=>X"0000001d0000001d0000001d0000001d", 10893=>X"0000001d0000001d0000001d0000001d", 10894=>X"0000001d0000001d0000001d0000001d", 
10895=>X"0000001d0000001d0000001d0000001d", 10896=>X"0000001d0000001d0000001d0000001d", 10897=>X"0000001d0000001d0000001d0000001d", 10898=>X"0000001d0000001d0000001d0000001d", 10899=>X"0000001d0000001d0000001d0000001d", 
10900=>X"0000001d0000001d0000001d0000001d", 10901=>X"0000001d0000001d0000001d0000001d", 10902=>X"0000001d0000001d0000001d0000001d", 10903=>X"0000001d0000001d0000001d0000001d", 10904=>X"0000001d0000001d0000001d0000001d", 
10905=>X"0000001d0000001d0000001d0000001d", 10906=>X"0000001d0000001d0000001d0000001d", 10907=>X"0000001d0000001d0000001d0000001d", 10908=>X"0000001d0000001d0000001d0000001d", 10909=>X"0000001d0000001d0000001d0000001d", 
10910=>X"0000001d0000001d0000001d0000001d", 10911=>X"0000001d0000001d0000001d0000001d", 10912=>X"0000001d0000001d0000001d0000001d", 10913=>X"0000001d0000001d0000001d0000001d", 10914=>X"0000001d0000001d0000001d0000001d", 
10915=>X"0000001d0000001d0000001d0000001d", 10916=>X"0000001d0000001d0000001d0000001d", 10917=>X"0000001d0000001d0000001d0000001d", 10918=>X"0000001d0000001d0000001d0000001d", 10919=>X"0000001d0000001d0000001d0000001d", 
10920=>X"0000001d0000001d0000001d0000001d", 10921=>X"0000001d0000001d0000001d0000001d", 10922=>X"0000001d0000001d0000001d0000001d", 10923=>X"0000001d0000001d0000001d0000001d", 10924=>X"0000001d0000001d0000001d0000001d", 
10925=>X"0000001d0000001d0000001d0000001d", 10926=>X"0000001d0000001d0000001d0000001d", 10927=>X"0000001d0000001d0000001d0000001d", 10928=>X"0000001d0000001d0000001d0000001d", 10929=>X"0000001d0000001d0000001d0000001d", 
10930=>X"0000001d0000001d0000001d0000001d", 10931=>X"0000001d0000001d0000001d0000001d", 10932=>X"0000001d0000001d0000001d0000001d", 10933=>X"0000001d0000001d0000001d0000001d", 10934=>X"0000001d0000001d0000001d0000001d", 
10935=>X"0000001d0000001d0000001d0000001d", 10936=>X"0000001d0000001d0000001d0000001d", 10937=>X"0000001d0000001d0000001d0000001d", 10938=>X"0000001d0000001d0000001d0000001d", 10939=>X"0000001d0000001d0000001d0000001d", 
10940=>X"0000001d0000001d0000001d0000001d", 10941=>X"0000001d0000001d0000001d0000001d", 10942=>X"0000001d0000001d0000001d0000001d", 10943=>X"0000001d0000001d0000001d0000001d", 10944=>X"0000001d0000001d0000001d0000001d", 
10945=>X"0000001d0000001d0000001d0000001d", 10946=>X"0000001d0000001d0000001d0000001d", 10947=>X"0000001d0000001d0000001d0000001d", 10948=>X"0000001d0000001d0000001d0000001d", 10949=>X"0000001d0000001d0000001d0000001d", 
10950=>X"0000001d0000001d0000001d0000001d", 10951=>X"0000001d0000001d0000001d0000001d", 10952=>X"0000001d0000001d0000001d0000001d", 10953=>X"0000001d0000001d0000001d0000001d", 10954=>X"0000001d0000001d0000001d0000001d", 
10955=>X"0000001d0000001d0000001d0000001d", 10956=>X"0000001d0000001d0000001d0000001d", 10957=>X"0000001d0000001d0000001d0000001d", 10958=>X"0000001d0000001d0000001d0000001d", 10959=>X"0000001d0000001d0000001d0000001d", 
10960=>X"0000001d0000001d0000001d0000001d", 10961=>X"0000001d0000001d0000001d0000001d", 10962=>X"0000001d0000001d0000001d0000001d", 10963=>X"0000001d0000001d0000001d0000001d", 10964=>X"0000001d0000001d0000001d0000001d", 
10965=>X"0000001d0000001d0000001d0000001d", 10966=>X"0000001d0000001d0000001d0000001d", 10967=>X"0000001d0000001d0000001d0000001d", 10968=>X"0000001d0000001d0000001d0000001d", 10969=>X"0000001d0000001d0000001d0000001d", 
10970=>X"0000001d0000001d0000001d0000001d", 10971=>X"0000001d0000001d0000001d0000001d", 10972=>X"0000001d0000001d0000001d0000001d", 10973=>X"0000001d0000001d0000001d0000001d", 10974=>X"0000001d0000001d0000001d0000001d", 
10975=>X"0000001d0000001d0000001d0000001d", 10976=>X"0000001d0000001d0000001d0000001d", 10977=>X"0000001d0000001d0000001d0000001d", 10978=>X"0000001d0000001d0000001d0000001d", 10979=>X"0000001d0000001d0000001d0000001d", 
10980=>X"0000001d0000001d0000001d0000001d", 10981=>X"0000001d0000001d0000001d0000001d", 10982=>X"0000001d0000001d0000001d0000001d", 10983=>X"0000001d0000001d0000001d0000001d", 10984=>X"0000001d0000001d0000001d0000001d", 
10985=>X"0000001d0000001d0000001d0000001d", 10986=>X"0000001d0000001d0000001d0000001d", 10987=>X"0000001d0000001d0000001d0000001d", 10988=>X"0000001d0000001d0000001d0000001d", 10989=>X"0000001d0000001d0000001d0000001d", 
10990=>X"0000001d0000001d0000001d0000001d", 10991=>X"0000001d0000001d0000001d0000001d", 10992=>X"0000001d0000001d0000001d0000001d", 10993=>X"0000001d0000001d0000001d0000001d", 10994=>X"0000001d0000001d0000001d0000001d", 
10995=>X"0000001d0000001d0000001d0000001d", 10996=>X"0000001d0000001d0000001d0000001d", 10997=>X"0000001d0000001d0000001d0000001d", 10998=>X"0000001d0000001d0000001d0000001d", 10999=>X"0000001d0000001d0000001d0000001d", 
11000=>X"0000001d0000001d0000001d0000001d", 11001=>X"0000001d0000001d0000001d0000001d", 11002=>X"0000001d0000001d0000001d0000001d", 11003=>X"0000001d0000001d0000001d0000001d", 11004=>X"0000001d0000001d0000001d0000001d", 
11005=>X"0000001d0000001d0000001d0000001d", 11006=>X"0000001d0000001d0000001d0000001d", 11007=>X"0000001d0000001d0000001d0000001d", 11008=>X"0000001d0000001d0000001d0000001d", 11009=>X"0000001d0000001d0000001d0000001d", 
11010=>X"0000001d0000001d0000001d0000001d", 11011=>X"0000001d0000001d0000001d0000001d", 11012=>X"0000001d0000001d0000001d0000001d", 11013=>X"0000001d0000001d0000001d0000001d", 11014=>X"0000001d0000001d0000001d0000001d", 
11015=>X"0000001d0000001d0000001d0000001d", 11016=>X"0000001d0000001d0000001d0000001d", 11017=>X"0000001d0000001d0000001d0000001d", 11018=>X"0000001d0000001d0000001d0000001d", 11019=>X"0000001d0000001d0000001d0000001d", 
11020=>X"0000001d0000001d0000001d0000001d", 11021=>X"0000001d0000001d0000001d0000001d", 11022=>X"0000001d0000001d0000001d0000001d", 11023=>X"0000001d0000001d0000001d0000001d", 11024=>X"0000001d0000001d0000001d0000001d", 
11025=>X"0000001d0000001d0000001d0000001d", 11026=>X"0000001d0000001d0000001d0000001d", 11027=>X"0000001d0000001d0000001d0000001d", 11028=>X"0000001d0000001d0000001d0000001d", 11029=>X"0000001d0000001d0000001d0000001d", 
11030=>X"0000001d0000001d0000001d0000001d", 11031=>X"0000001d0000001d0000001d0000001d", 11032=>X"0000001d0000001d0000001d0000001d", 11033=>X"0000001d0000001d0000001d0000001d", 11034=>X"0000001d0000001d0000001d0000001d", 
11035=>X"0000001d0000001d0000001d0000001d", 11036=>X"0000001d0000001d0000001d0000001d", 11037=>X"0000001d0000001d0000001d0000001d", 11038=>X"0000001d0000001d0000001d0000001d", 11039=>X"0000001d0000001d0000001d0000001d", 
11040=>X"0000001d0000001d0000001d0000001d", 11041=>X"0000001d0000001d0000001d0000001d", 11042=>X"0000001d0000001d0000001d0000001d", 11043=>X"0000001d0000001d0000001d0000001d", 11044=>X"0000001d0000001d0000001d0000001d", 
11045=>X"0000001d0000001d0000001d0000001d", 11046=>X"0000001d0000001d0000001d0000001d", 11047=>X"0000001d0000001d0000001d0000001d", 11048=>X"0000001d0000001d0000001d0000001d", 11049=>X"0000001d0000001d0000001d0000001d", 
11050=>X"0000001d0000001d0000001d0000001d", 11051=>X"0000001d0000001d0000001d0000001d", 11052=>X"0000001d0000001d0000001d0000001d", 11053=>X"0000001d0000001d0000001d0000001d", 11054=>X"0000001d0000001d0000001d0000001d", 
11055=>X"0000001d0000001d0000001d0000001d", 11056=>X"0000001d0000001d0000001d0000001d", 11057=>X"0000001d0000001d0000001d0000001d", 11058=>X"0000001d0000001d0000001d0000001d", 11059=>X"0000001d0000001d0000001d0000001d", 
11060=>X"0000001d0000001d0000001d0000001d", 11061=>X"0000001d0000001d0000001d0000001d", 11062=>X"0000001d0000001d0000001d0000001d", 11063=>X"0000001d0000001d0000001d0000001d", 11064=>X"0000001d0000001d0000001d0000001d", 
11065=>X"0000001d0000001d0000001d0000001d", 11066=>X"0000001d0000001d0000001d0000001d", 11067=>X"0000001d0000001d0000001d0000001d", 11068=>X"0000001c0000001c0000001c0000001c", 11069=>X"0000001c0000001c0000001c0000001c", 
11070=>X"0000001c0000001c0000001c0000001c", 11071=>X"0000001c0000001c0000001c0000001c", 11072=>X"0000001c0000001c0000001c0000001c", 11073=>X"0000001c0000001c0000001c0000001c", 11074=>X"0000001c0000001c0000001c0000001c", 
11075=>X"0000001c0000001c0000001c0000001c", 11076=>X"0000001c0000001c0000001c0000001c", 11077=>X"0000001c0000001c0000001c0000001c", 11078=>X"0000001c0000001c0000001c0000001c", 11079=>X"0000001c0000001c0000001c0000001c", 
11080=>X"0000001c0000001c0000001c0000001c", 11081=>X"0000001c0000001c0000001c0000001c", 11082=>X"0000001c0000001c0000001c0000001c", 11083=>X"0000001c0000001c0000001c0000001c", 11084=>X"0000001c0000001c0000001c0000001c", 
11085=>X"0000001c0000001c0000001c0000001c", 11086=>X"0000001c0000001c0000001c0000001c", 11087=>X"0000001c0000001c0000001c0000001c", 11088=>X"0000001c0000001c0000001c0000001c", 11089=>X"0000001c0000001c0000001c0000001c", 
11090=>X"0000001c0000001c0000001c0000001c", 11091=>X"0000001c0000001c0000001c0000001c", 11092=>X"0000001c0000001c0000001c0000001c", 11093=>X"0000001c0000001c0000001c0000001c", 11094=>X"0000001c0000001c0000001c0000001c", 
11095=>X"0000001c0000001c0000001c0000001c", 11096=>X"0000001c0000001c0000001c0000001c", 11097=>X"0000001c0000001c0000001c0000001c", 11098=>X"0000001c0000001c0000001c0000001c", 11099=>X"0000001c0000001c0000001c0000001c", 
11100=>X"0000001c0000001c0000001c0000001c", 11101=>X"0000001c0000001c0000001c0000001c", 11102=>X"0000001c0000001c0000001c0000001c", 11103=>X"0000001c0000001c0000001c0000001c", 11104=>X"0000001c0000001c0000001c0000001c", 
11105=>X"0000001c0000001c0000001c0000001c", 11106=>X"0000001c0000001c0000001c0000001c", 11107=>X"0000001c0000001c0000001c0000001c", 11108=>X"0000001c0000001c0000001c0000001c", 11109=>X"0000001c0000001c0000001c0000001c", 
11110=>X"0000001c0000001c0000001c0000001c", 11111=>X"0000001c0000001c0000001c0000001c", 11112=>X"0000001c0000001c0000001c0000001c", 11113=>X"0000001c0000001c0000001c0000001c", 11114=>X"0000001c0000001c0000001c0000001c", 
11115=>X"0000001c0000001c0000001c0000001c", 11116=>X"0000001c0000001c0000001c0000001c", 11117=>X"0000001c0000001c0000001c0000001c", 11118=>X"0000001c0000001c0000001c0000001c", 11119=>X"0000001c0000001c0000001c0000001c", 
11120=>X"0000001c0000001c0000001c0000001c", 11121=>X"0000001c0000001c0000001c0000001c", 11122=>X"0000001c0000001c0000001c0000001c", 11123=>X"0000001c0000001c0000001c0000001c", 11124=>X"0000001c0000001c0000001c0000001c", 
11125=>X"0000001c0000001c0000001c0000001c", 11126=>X"0000001c0000001c0000001c0000001c", 11127=>X"0000001c0000001c0000001c0000001c", 11128=>X"0000001c0000001c0000001c0000001c", 11129=>X"0000001c0000001c0000001c0000001c", 
11130=>X"0000001c0000001c0000001c0000001c", 11131=>X"0000001c0000001c0000001c0000001c", 11132=>X"0000001c0000001c0000001c0000001c", 11133=>X"0000001c0000001c0000001c0000001c", 11134=>X"0000001c0000001c0000001c0000001c", 
11135=>X"0000001c0000001c0000001c0000001c", 11136=>X"0000001c0000001c0000001c0000001c", 11137=>X"0000001c0000001c0000001c0000001c", 11138=>X"0000001c0000001c0000001c0000001c", 11139=>X"0000001c0000001c0000001c0000001c", 
11140=>X"0000001c0000001c0000001c0000001c", 11141=>X"0000001c0000001c0000001c0000001c", 11142=>X"0000001c0000001c0000001c0000001c", 11143=>X"0000001c0000001c0000001c0000001c", 11144=>X"0000001c0000001c0000001c0000001c", 
11145=>X"0000001c0000001c0000001c0000001c", 11146=>X"0000001c0000001c0000001c0000001c", 11147=>X"0000001c0000001c0000001c0000001c", 11148=>X"0000001c0000001c0000001c0000001c", 11149=>X"0000001c0000001c0000001c0000001c", 
11150=>X"0000001c0000001c0000001c0000001c", 11151=>X"0000001c0000001c0000001c0000001c", 11152=>X"0000001c0000001c0000001c0000001c", 11153=>X"0000001c0000001c0000001c0000001c", 11154=>X"0000001c0000001c0000001c0000001c", 
11155=>X"0000001c0000001c0000001c0000001c", 11156=>X"0000001c0000001c0000001c0000001c", 11157=>X"0000001c0000001c0000001c0000001c", 11158=>X"0000001c0000001c0000001c0000001c", 11159=>X"0000001c0000001c0000001c0000001c", 
11160=>X"0000001c0000001c0000001c0000001c", 11161=>X"0000001c0000001c0000001c0000001c", 11162=>X"0000001c0000001c0000001c0000001c", 11163=>X"0000001c0000001c0000001c0000001c", 11164=>X"0000001c0000001c0000001c0000001c", 
11165=>X"0000001c0000001c0000001c0000001c", 11166=>X"0000001c0000001c0000001c0000001c", 11167=>X"0000001c0000001c0000001c0000001c", 11168=>X"0000001c0000001c0000001c0000001c", 11169=>X"0000001c0000001c0000001c0000001c", 
11170=>X"0000001c0000001c0000001c0000001c", 11171=>X"0000001c0000001c0000001c0000001c", 11172=>X"0000001c0000001c0000001c0000001c", 11173=>X"0000001c0000001c0000001c0000001c", 11174=>X"0000001c0000001c0000001c0000001c", 
11175=>X"0000001c0000001c0000001c0000001c", 11176=>X"0000001c0000001c0000001c0000001c", 11177=>X"0000001c0000001c0000001c0000001c", 11178=>X"0000001c0000001c0000001c0000001c", 11179=>X"0000001c0000001c0000001c0000001c", 
11180=>X"0000001c0000001c0000001c0000001c", 11181=>X"0000001c0000001c0000001c0000001c", 11182=>X"0000001c0000001c0000001c0000001c", 11183=>X"0000001c0000001c0000001c0000001c", 11184=>X"0000001c0000001c0000001c0000001c", 
11185=>X"0000001c0000001c0000001c0000001c", 11186=>X"0000001c0000001c0000001c0000001c", 11187=>X"0000001c0000001c0000001c0000001c", 11188=>X"0000001c0000001c0000001c0000001c", 11189=>X"0000001c0000001c0000001c0000001c", 
11190=>X"0000001c0000001c0000001c0000001c", 11191=>X"0000001c0000001c0000001c0000001c", 11192=>X"0000001c0000001c0000001c0000001c", 11193=>X"0000001c0000001c0000001c0000001c", 11194=>X"0000001c0000001c0000001c0000001c", 
11195=>X"0000001c0000001c0000001c0000001c", 11196=>X"0000001c0000001c0000001c0000001c", 11197=>X"0000001c0000001c0000001c0000001c", 11198=>X"0000001c0000001c0000001c0000001c", 11199=>X"0000001c0000001c0000001c0000001c", 
11200=>X"0000001c0000001c0000001c0000001c", 11201=>X"0000001c0000001c0000001c0000001c", 11202=>X"0000001c0000001c0000001c0000001c", 11203=>X"0000001c0000001c0000001c0000001c", 11204=>X"0000001c0000001c0000001c0000001c", 
11205=>X"0000001c0000001c0000001c0000001c", 11206=>X"0000001c0000001c0000001c0000001c", 11207=>X"0000001c0000001c0000001c0000001c", 11208=>X"0000001c0000001c0000001c0000001c", 11209=>X"0000001c0000001c0000001c0000001c", 
11210=>X"0000001c0000001c0000001c0000001c", 11211=>X"0000001c0000001c0000001c0000001c", 11212=>X"0000001c0000001c0000001c0000001c", 11213=>X"0000001c0000001c0000001c0000001c", 11214=>X"0000001c0000001c0000001c0000001c", 
11215=>X"0000001c0000001c0000001c0000001c", 11216=>X"0000001c0000001c0000001c0000001c", 11217=>X"0000001c0000001c0000001c0000001c", 11218=>X"0000001c0000001c0000001c0000001c", 11219=>X"0000001c0000001c0000001c0000001c", 
11220=>X"0000001c0000001c0000001c0000001c", 11221=>X"0000001c0000001c0000001c0000001c", 11222=>X"0000001c0000001c0000001c0000001c", 11223=>X"0000001c0000001c0000001c0000001c", 11224=>X"0000001c0000001c0000001c0000001c", 
11225=>X"0000001c0000001c0000001c0000001c", 11226=>X"0000001c0000001c0000001c0000001c", 11227=>X"0000001c0000001c0000001c0000001c", 11228=>X"0000001c0000001c0000001c0000001c", 11229=>X"0000001c0000001c0000001c0000001c", 
11230=>X"0000001c0000001c0000001c0000001c", 11231=>X"0000001c0000001c0000001c0000001c", 11232=>X"0000001c0000001c0000001c0000001c", 11233=>X"0000001c0000001c0000001c0000001c", 11234=>X"0000001c0000001c0000001c0000001c", 
11235=>X"0000001c0000001c0000001c0000001c", 11236=>X"0000001c0000001c0000001c0000001c", 11237=>X"0000001c0000001c0000001c0000001c", 11238=>X"0000001c0000001c0000001c0000001c", 11239=>X"0000001c0000001c0000001c0000001c", 
11240=>X"0000001c0000001c0000001c0000001c", 11241=>X"0000001c0000001c0000001c0000001c", 11242=>X"0000001c0000001c0000001c0000001c", 11243=>X"0000001c0000001c0000001c0000001c", 11244=>X"0000001c0000001c0000001c0000001c", 
11245=>X"0000001c0000001c0000001c0000001c", 11246=>X"0000001c0000001c0000001c0000001c", 11247=>X"0000001c0000001c0000001c0000001c", 11248=>X"0000001c0000001c0000001c0000001c", 11249=>X"0000001c0000001c0000001c0000001c", 
11250=>X"0000001c0000001c0000001c0000001c", 11251=>X"0000001c0000001c0000001c0000001c", 11252=>X"0000001c0000001c0000001c0000001c", 11253=>X"0000001c0000001c0000001c0000001c", 11254=>X"0000001c0000001c0000001c0000001c", 
11255=>X"0000001c0000001c0000001c0000001c", 11256=>X"0000001c0000001c0000001c0000001c", 11257=>X"0000001c0000001c0000001c0000001c", 11258=>X"0000001c0000001c0000001c0000001c", 11259=>X"0000001c0000001c0000001c0000001c", 
11260=>X"0000001c0000001c0000001c0000001c", 11261=>X"0000001c0000001c0000001c0000001c", 11262=>X"0000001c0000001c0000001c0000001c", 11263=>X"0000001c0000001c0000001c0000001c", 11264=>X"0000001c0000001c0000001c0000001c", 
11265=>X"0000001c0000001c0000001c0000001c", 11266=>X"0000001c0000001c0000001c0000001c", 11267=>X"0000001c0000001c0000001c0000001c", 11268=>X"0000001c0000001c0000001c0000001c", 11269=>X"0000001c0000001c0000001c0000001c", 
11270=>X"0000001c0000001c0000001c0000001c", 11271=>X"0000001c0000001c0000001c0000001c", 11272=>X"0000001c0000001c0000001c0000001c", 11273=>X"0000001c0000001c0000001c0000001c", 11274=>X"0000001c0000001c0000001c0000001c", 
11275=>X"0000001c0000001c0000001c0000001c", 11276=>X"0000001c0000001c0000001c0000001c", 11277=>X"0000001c0000001c0000001c0000001c", 11278=>X"0000001c0000001c0000001c0000001c", 11279=>X"0000001c0000001c0000001c0000001c", 
11280=>X"0000001c0000001c0000001c0000001c", 11281=>X"0000001c0000001c0000001c0000001c", 11282=>X"0000001c0000001c0000001c0000001c", 11283=>X"0000001c0000001c0000001c0000001c", 11284=>X"0000001c0000001c0000001c0000001c", 
11285=>X"0000001c0000001c0000001c0000001c", 11286=>X"0000001c0000001c0000001c0000001c", 11287=>X"0000001c0000001c0000001c0000001c", 11288=>X"0000001c0000001c0000001c0000001c", 11289=>X"0000001c0000001c0000001c0000001c", 
11290=>X"0000001c0000001c0000001c0000001c", 11291=>X"0000001c0000001c0000001c0000001c", 11292=>X"0000001c0000001c0000001c0000001c", 11293=>X"0000001c0000001c0000001c0000001c", 11294=>X"0000001c0000001c0000001c0000001c", 
11295=>X"0000001c0000001c0000001c0000001c", 11296=>X"0000001c0000001c0000001c0000001c", 11297=>X"0000001c0000001c0000001c0000001c", 11298=>X"0000001c0000001c0000001c0000001c", 11299=>X"0000001c0000001c0000001c0000001c", 
11300=>X"0000001c0000001c0000001c0000001c", 11301=>X"0000001c0000001c0000001c0000001c", 11302=>X"0000001c0000001c0000001c0000001c", 11303=>X"0000001c0000001c0000001c0000001c", 11304=>X"0000001c0000001c0000001c0000001c", 
11305=>X"0000001c0000001c0000001c0000001c", 11306=>X"0000001c0000001c0000001c0000001c", 11307=>X"0000001c0000001c0000001c0000001c", 11308=>X"0000001c0000001c0000001c0000001c", 11309=>X"0000001c0000001c0000001c0000001c", 
11310=>X"0000001c0000001c0000001c0000001c", 11311=>X"0000001c0000001c0000001c0000001c", 11312=>X"0000001c0000001c0000001c0000001c", 11313=>X"0000001c0000001c0000001c0000001c", 11314=>X"0000001c0000001c0000001c0000001c", 
11315=>X"0000001c0000001c0000001c0000001c", 11316=>X"0000001c0000001c0000001c0000001c", 11317=>X"0000001c0000001c0000001c0000001c", 11318=>X"0000001c0000001c0000001c0000001c", 11319=>X"0000001c0000001c0000001c0000001c", 
11320=>X"0000001c0000001c0000001c0000001c", 11321=>X"0000001c0000001c0000001c0000001c", 11322=>X"0000001c0000001c0000001c0000001c", 11323=>X"0000001c0000001c0000001c0000001c", 11324=>X"0000001c0000001c0000001c0000001c", 
11325=>X"0000001c0000001c0000001c0000001c", 11326=>X"0000001c0000001c0000001c0000001c", 11327=>X"0000001c0000001c0000001c0000001c", 11328=>X"0000001c0000001c0000001c0000001c", 11329=>X"0000001c0000001c0000001c0000001c", 
11330=>X"0000001c0000001c0000001c0000001c", 11331=>X"0000001c0000001c0000001c0000001c", 11332=>X"0000001c0000001c0000001c0000001c", 11333=>X"0000001c0000001c0000001c0000001c", 11334=>X"0000001c0000001c0000001c0000001c", 
11335=>X"0000001c0000001c0000001c0000001c", 11336=>X"0000001c0000001c0000001c0000001c", 11337=>X"0000001c0000001c0000001c0000001c", 11338=>X"0000001c0000001c0000001c0000001c", 11339=>X"0000001c0000001c0000001c0000001c", 
11340=>X"0000001c0000001c0000001c0000001c", 11341=>X"0000001c0000001c0000001c0000001c", 11342=>X"0000001c0000001c0000001c0000001c", 11343=>X"0000001c0000001c0000001c0000001c", 11344=>X"0000001c0000001c0000001c0000001c", 
11345=>X"0000001c0000001c0000001c0000001c", 11346=>X"0000001c0000001c0000001c0000001c", 11347=>X"0000001c0000001c0000001c0000001c", 11348=>X"0000001c0000001c0000001c0000001c", 11349=>X"0000001c0000001c0000001c0000001c", 
11350=>X"0000001c0000001c0000001c0000001c", 11351=>X"0000001c0000001c0000001c0000001c", 11352=>X"0000001c0000001c0000001c0000001c", 11353=>X"0000001c0000001c0000001c0000001c", 11354=>X"0000001c0000001c0000001c0000001c", 
11355=>X"0000001c0000001c0000001c0000001c", 11356=>X"0000001c0000001c0000001c0000001c", 11357=>X"0000001c0000001c0000001c0000001c", 11358=>X"0000001c0000001c0000001c0000001c", 11359=>X"0000001c0000001c0000001c0000001c", 
11360=>X"0000001c0000001c0000001c0000001c", 11361=>X"0000001c0000001c0000001c0000001c", 11362=>X"0000001c0000001c0000001c0000001c", 11363=>X"0000001c0000001c0000001c0000001c", 11364=>X"0000001c0000001c0000001c0000001c", 
11365=>X"0000001c0000001c0000001c0000001c", 11366=>X"0000001c0000001c0000001c0000001c", 11367=>X"0000001c0000001c0000001c0000001c", 11368=>X"0000001c0000001c0000001c0000001c", 11369=>X"0000001c0000001c0000001c0000001c", 
11370=>X"0000001c0000001c0000001c0000001c", 11371=>X"0000001c0000001c0000001c0000001c", 11372=>X"0000001c0000001c0000001c0000001c", 11373=>X"0000001c0000001c0000001c0000001c", 11374=>X"0000001c0000001c0000001c0000001c", 
11375=>X"0000001c0000001c0000001c0000001c", 11376=>X"0000001c0000001c0000001c0000001c", 11377=>X"0000001c0000001c0000001c0000001c", 11378=>X"0000001c0000001c0000001c0000001c", 11379=>X"0000001c0000001c0000001c0000001c", 
11380=>X"0000001c0000001c0000001c0000001c", 11381=>X"0000001c0000001c0000001c0000001c", 11382=>X"0000001c0000001c0000001c0000001c", 11383=>X"0000001c0000001c0000001c0000001c", 11384=>X"0000001c0000001c0000001c0000001c", 
11385=>X"0000001c0000001c0000001c0000001c", 11386=>X"0000001c0000001c0000001c0000001c", 11387=>X"0000001c0000001c0000001c0000001c", 11388=>X"0000001c0000001c0000001c0000001c", 11389=>X"0000001c0000001c0000001c0000001c", 
11390=>X"0000001c0000001c0000001c0000001c", 11391=>X"0000001c0000001c0000001c0000001c", 11392=>X"0000001c0000001c0000001c0000001c", 11393=>X"0000001c0000001c0000001c0000001c", 11394=>X"0000001c0000001c0000001c0000001c", 
11395=>X"0000001c0000001c0000001c0000001c", 11396=>X"0000001c0000001c0000001c0000001c", 11397=>X"0000001c0000001c0000001c0000001c", 11398=>X"0000001c0000001c0000001c0000001c", 11399=>X"0000001c0000001c0000001c0000001c", 
11400=>X"0000001c0000001c0000001c0000001c", 11401=>X"0000001c0000001c0000001c0000001c", 11402=>X"0000001b0000001b0000001c0000001c", 11403=>X"0000001b0000001b0000001b0000001b", 11404=>X"0000001b0000001b0000001b0000001b", 
11405=>X"0000001b0000001b0000001b0000001b", 11406=>X"0000001b0000001b0000001b0000001b", 11407=>X"0000001b0000001b0000001b0000001b", 11408=>X"0000001b0000001b0000001b0000001b", 11409=>X"0000001b0000001b0000001b0000001b", 
11410=>X"0000001b0000001b0000001b0000001b", 11411=>X"0000001b0000001b0000001b0000001b", 11412=>X"0000001b0000001b0000001b0000001b", 11413=>X"0000001b0000001b0000001b0000001b", 11414=>X"0000001b0000001b0000001b0000001b", 
11415=>X"0000001b0000001b0000001b0000001b", 11416=>X"0000001b0000001b0000001b0000001b", 11417=>X"0000001b0000001b0000001b0000001b", 11418=>X"0000001b0000001b0000001b0000001b", 11419=>X"0000001b0000001b0000001b0000001b", 
11420=>X"0000001b0000001b0000001b0000001b", 11421=>X"0000001b0000001b0000001b0000001b", 11422=>X"0000001b0000001b0000001b0000001b", 11423=>X"0000001b0000001b0000001b0000001b", 11424=>X"0000001b0000001b0000001b0000001b", 
11425=>X"0000001b0000001b0000001b0000001b", 11426=>X"0000001b0000001b0000001b0000001b", 11427=>X"0000001b0000001b0000001b0000001b", 11428=>X"0000001b0000001b0000001b0000001b", 11429=>X"0000001b0000001b0000001b0000001b", 
11430=>X"0000001b0000001b0000001b0000001b", 11431=>X"0000001b0000001b0000001b0000001b", 11432=>X"0000001b0000001b0000001b0000001b", 11433=>X"0000001b0000001b0000001b0000001b", 11434=>X"0000001b0000001b0000001b0000001b", 
11435=>X"0000001b0000001b0000001b0000001b", 11436=>X"0000001b0000001b0000001b0000001b", 11437=>X"0000001b0000001b0000001b0000001b", 11438=>X"0000001b0000001b0000001b0000001b", 11439=>X"0000001b0000001b0000001b0000001b", 
11440=>X"0000001b0000001b0000001b0000001b", 11441=>X"0000001b0000001b0000001b0000001b", 11442=>X"0000001b0000001b0000001b0000001b", 11443=>X"0000001b0000001b0000001b0000001b", 11444=>X"0000001b0000001b0000001b0000001b", 
11445=>X"0000001b0000001b0000001b0000001b", 11446=>X"0000001b0000001b0000001b0000001b", 11447=>X"0000001b0000001b0000001b0000001b", 11448=>X"0000001b0000001b0000001b0000001b", 11449=>X"0000001b0000001b0000001b0000001b", 
11450=>X"0000001b0000001b0000001b0000001b", 11451=>X"0000001b0000001b0000001b0000001b", 11452=>X"0000001b0000001b0000001b0000001b", 11453=>X"0000001b0000001b0000001b0000001b", 11454=>X"0000001b0000001b0000001b0000001b", 
11455=>X"0000001b0000001b0000001b0000001b", 11456=>X"0000001b0000001b0000001b0000001b", 11457=>X"0000001b0000001b0000001b0000001b", 11458=>X"0000001b0000001b0000001b0000001b", 11459=>X"0000001b0000001b0000001b0000001b", 
11460=>X"0000001b0000001b0000001b0000001b", 11461=>X"0000001b0000001b0000001b0000001b", 11462=>X"0000001b0000001b0000001b0000001b", 11463=>X"0000001b0000001b0000001b0000001b", 11464=>X"0000001b0000001b0000001b0000001b", 
11465=>X"0000001b0000001b0000001b0000001b", 11466=>X"0000001b0000001b0000001b0000001b", 11467=>X"0000001b0000001b0000001b0000001b", 11468=>X"0000001b0000001b0000001b0000001b", 11469=>X"0000001b0000001b0000001b0000001b", 
11470=>X"0000001b0000001b0000001b0000001b", 11471=>X"0000001b0000001b0000001b0000001b", 11472=>X"0000001b0000001b0000001b0000001b", 11473=>X"0000001b0000001b0000001b0000001b", 11474=>X"0000001b0000001b0000001b0000001b", 
11475=>X"0000001b0000001b0000001b0000001b", 11476=>X"0000001b0000001b0000001b0000001b", 11477=>X"0000001b0000001b0000001b0000001b", 11478=>X"0000001b0000001b0000001b0000001b", 11479=>X"0000001b0000001b0000001b0000001b", 
11480=>X"0000001b0000001b0000001b0000001b", 11481=>X"0000001b0000001b0000001b0000001b", 11482=>X"0000001b0000001b0000001b0000001b", 11483=>X"0000001b0000001b0000001b0000001b", 11484=>X"0000001b0000001b0000001b0000001b", 
11485=>X"0000001b0000001b0000001b0000001b", 11486=>X"0000001b0000001b0000001b0000001b", 11487=>X"0000001b0000001b0000001b0000001b", 11488=>X"0000001b0000001b0000001b0000001b", 11489=>X"0000001b0000001b0000001b0000001b", 
11490=>X"0000001b0000001b0000001b0000001b", 11491=>X"0000001b0000001b0000001b0000001b", 11492=>X"0000001b0000001b0000001b0000001b", 11493=>X"0000001b0000001b0000001b0000001b", 11494=>X"0000001b0000001b0000001b0000001b", 
11495=>X"0000001b0000001b0000001b0000001b", 11496=>X"0000001b0000001b0000001b0000001b", 11497=>X"0000001b0000001b0000001b0000001b", 11498=>X"0000001b0000001b0000001b0000001b", 11499=>X"0000001b0000001b0000001b0000001b", 
11500=>X"0000001b0000001b0000001b0000001b", 11501=>X"0000001b0000001b0000001b0000001b", 11502=>X"0000001b0000001b0000001b0000001b", 11503=>X"0000001b0000001b0000001b0000001b", 11504=>X"0000001b0000001b0000001b0000001b", 
11505=>X"0000001b0000001b0000001b0000001b", 11506=>X"0000001b0000001b0000001b0000001b", 11507=>X"0000001b0000001b0000001b0000001b", 11508=>X"0000001b0000001b0000001b0000001b", 11509=>X"0000001b0000001b0000001b0000001b", 
11510=>X"0000001b0000001b0000001b0000001b", 11511=>X"0000001b0000001b0000001b0000001b", 11512=>X"0000001b0000001b0000001b0000001b", 11513=>X"0000001b0000001b0000001b0000001b", 11514=>X"0000001b0000001b0000001b0000001b", 
11515=>X"0000001b0000001b0000001b0000001b", 11516=>X"0000001b0000001b0000001b0000001b", 11517=>X"0000001b0000001b0000001b0000001b", 11518=>X"0000001b0000001b0000001b0000001b", 11519=>X"0000001b0000001b0000001b0000001b", 
11520=>X"0000001b0000001b0000001b0000001b", 11521=>X"0000001b0000001b0000001b0000001b", 11522=>X"0000001b0000001b0000001b0000001b", 11523=>X"0000001b0000001b0000001b0000001b", 11524=>X"0000001b0000001b0000001b0000001b", 
11525=>X"0000001b0000001b0000001b0000001b", 11526=>X"0000001b0000001b0000001b0000001b", 11527=>X"0000001b0000001b0000001b0000001b", 11528=>X"0000001b0000001b0000001b0000001b", 11529=>X"0000001b0000001b0000001b0000001b", 
11530=>X"0000001b0000001b0000001b0000001b", 11531=>X"0000001b0000001b0000001b0000001b", 11532=>X"0000001b0000001b0000001b0000001b", 11533=>X"0000001b0000001b0000001b0000001b", 11534=>X"0000001b0000001b0000001b0000001b", 
11535=>X"0000001b0000001b0000001b0000001b", 11536=>X"0000001b0000001b0000001b0000001b", 11537=>X"0000001b0000001b0000001b0000001b", 11538=>X"0000001b0000001b0000001b0000001b", 11539=>X"0000001b0000001b0000001b0000001b", 
11540=>X"0000001b0000001b0000001b0000001b", 11541=>X"0000001b0000001b0000001b0000001b", 11542=>X"0000001b0000001b0000001b0000001b", 11543=>X"0000001b0000001b0000001b0000001b", 11544=>X"0000001b0000001b0000001b0000001b", 
11545=>X"0000001b0000001b0000001b0000001b", 11546=>X"0000001b0000001b0000001b0000001b", 11547=>X"0000001b0000001b0000001b0000001b", 11548=>X"0000001b0000001b0000001b0000001b", 11549=>X"0000001b0000001b0000001b0000001b", 
11550=>X"0000001b0000001b0000001b0000001b", 11551=>X"0000001b0000001b0000001b0000001b", 11552=>X"0000001b0000001b0000001b0000001b", 11553=>X"0000001b0000001b0000001b0000001b", 11554=>X"0000001b0000001b0000001b0000001b", 
11555=>X"0000001b0000001b0000001b0000001b", 11556=>X"0000001b0000001b0000001b0000001b", 11557=>X"0000001b0000001b0000001b0000001b", 11558=>X"0000001b0000001b0000001b0000001b", 11559=>X"0000001b0000001b0000001b0000001b", 
11560=>X"0000001b0000001b0000001b0000001b", 11561=>X"0000001b0000001b0000001b0000001b", 11562=>X"0000001b0000001b0000001b0000001b", 11563=>X"0000001b0000001b0000001b0000001b", 11564=>X"0000001b0000001b0000001b0000001b", 
11565=>X"0000001b0000001b0000001b0000001b", 11566=>X"0000001b0000001b0000001b0000001b", 11567=>X"0000001b0000001b0000001b0000001b", 11568=>X"0000001b0000001b0000001b0000001b", 11569=>X"0000001b0000001b0000001b0000001b", 
11570=>X"0000001b0000001b0000001b0000001b", 11571=>X"0000001b0000001b0000001b0000001b", 11572=>X"0000001b0000001b0000001b0000001b", 11573=>X"0000001b0000001b0000001b0000001b", 11574=>X"0000001b0000001b0000001b0000001b", 
11575=>X"0000001b0000001b0000001b0000001b", 11576=>X"0000001b0000001b0000001b0000001b", 11577=>X"0000001b0000001b0000001b0000001b", 11578=>X"0000001b0000001b0000001b0000001b", 11579=>X"0000001b0000001b0000001b0000001b", 
11580=>X"0000001b0000001b0000001b0000001b", 11581=>X"0000001b0000001b0000001b0000001b", 11582=>X"0000001b0000001b0000001b0000001b", 11583=>X"0000001b0000001b0000001b0000001b", 11584=>X"0000001b0000001b0000001b0000001b", 
11585=>X"0000001b0000001b0000001b0000001b", 11586=>X"0000001b0000001b0000001b0000001b", 11587=>X"0000001b0000001b0000001b0000001b", 11588=>X"0000001b0000001b0000001b0000001b", 11589=>X"0000001b0000001b0000001b0000001b", 
11590=>X"0000001b0000001b0000001b0000001b", 11591=>X"0000001b0000001b0000001b0000001b", 11592=>X"0000001b0000001b0000001b0000001b", 11593=>X"0000001b0000001b0000001b0000001b", 11594=>X"0000001b0000001b0000001b0000001b", 
11595=>X"0000001b0000001b0000001b0000001b", 11596=>X"0000001b0000001b0000001b0000001b", 11597=>X"0000001b0000001b0000001b0000001b", 11598=>X"0000001b0000001b0000001b0000001b", 11599=>X"0000001b0000001b0000001b0000001b", 
11600=>X"0000001b0000001b0000001b0000001b", 11601=>X"0000001b0000001b0000001b0000001b", 11602=>X"0000001b0000001b0000001b0000001b", 11603=>X"0000001b0000001b0000001b0000001b", 11604=>X"0000001b0000001b0000001b0000001b", 
11605=>X"0000001b0000001b0000001b0000001b", 11606=>X"0000001b0000001b0000001b0000001b", 11607=>X"0000001b0000001b0000001b0000001b", 11608=>X"0000001b0000001b0000001b0000001b", 11609=>X"0000001b0000001b0000001b0000001b", 
11610=>X"0000001b0000001b0000001b0000001b", 11611=>X"0000001b0000001b0000001b0000001b", 11612=>X"0000001b0000001b0000001b0000001b", 11613=>X"0000001b0000001b0000001b0000001b", 11614=>X"0000001b0000001b0000001b0000001b", 
11615=>X"0000001b0000001b0000001b0000001b", 11616=>X"0000001b0000001b0000001b0000001b", 11617=>X"0000001b0000001b0000001b0000001b", 11618=>X"0000001b0000001b0000001b0000001b", 11619=>X"0000001b0000001b0000001b0000001b", 
11620=>X"0000001b0000001b0000001b0000001b", 11621=>X"0000001b0000001b0000001b0000001b", 11622=>X"0000001b0000001b0000001b0000001b", 11623=>X"0000001b0000001b0000001b0000001b", 11624=>X"0000001b0000001b0000001b0000001b", 
11625=>X"0000001b0000001b0000001b0000001b", 11626=>X"0000001b0000001b0000001b0000001b", 11627=>X"0000001b0000001b0000001b0000001b", 11628=>X"0000001b0000001b0000001b0000001b", 11629=>X"0000001b0000001b0000001b0000001b", 
11630=>X"0000001b0000001b0000001b0000001b", 11631=>X"0000001b0000001b0000001b0000001b", 11632=>X"0000001b0000001b0000001b0000001b", 11633=>X"0000001b0000001b0000001b0000001b", 11634=>X"0000001b0000001b0000001b0000001b", 
11635=>X"0000001b0000001b0000001b0000001b", 11636=>X"0000001b0000001b0000001b0000001b", 11637=>X"0000001b0000001b0000001b0000001b", 11638=>X"0000001b0000001b0000001b0000001b", 11639=>X"0000001b0000001b0000001b0000001b", 
11640=>X"0000001b0000001b0000001b0000001b", 11641=>X"0000001b0000001b0000001b0000001b", 11642=>X"0000001b0000001b0000001b0000001b", 11643=>X"0000001b0000001b0000001b0000001b", 11644=>X"0000001b0000001b0000001b0000001b", 
11645=>X"0000001b0000001b0000001b0000001b", 11646=>X"0000001b0000001b0000001b0000001b", 11647=>X"0000001b0000001b0000001b0000001b", 11648=>X"0000001b0000001b0000001b0000001b", 11649=>X"0000001b0000001b0000001b0000001b", 
11650=>X"0000001b0000001b0000001b0000001b", 11651=>X"0000001b0000001b0000001b0000001b", 11652=>X"0000001b0000001b0000001b0000001b", 11653=>X"0000001b0000001b0000001b0000001b", 11654=>X"0000001b0000001b0000001b0000001b", 
11655=>X"0000001b0000001b0000001b0000001b", 11656=>X"0000001b0000001b0000001b0000001b", 11657=>X"0000001b0000001b0000001b0000001b", 11658=>X"0000001b0000001b0000001b0000001b", 11659=>X"0000001b0000001b0000001b0000001b", 
11660=>X"0000001b0000001b0000001b0000001b", 11661=>X"0000001b0000001b0000001b0000001b", 11662=>X"0000001b0000001b0000001b0000001b", 11663=>X"0000001b0000001b0000001b0000001b", 11664=>X"0000001b0000001b0000001b0000001b", 
11665=>X"0000001b0000001b0000001b0000001b", 11666=>X"0000001b0000001b0000001b0000001b", 11667=>X"0000001b0000001b0000001b0000001b", 11668=>X"0000001b0000001b0000001b0000001b", 11669=>X"0000001b0000001b0000001b0000001b", 
11670=>X"0000001b0000001b0000001b0000001b", 11671=>X"0000001b0000001b0000001b0000001b", 11672=>X"0000001b0000001b0000001b0000001b", 11673=>X"0000001b0000001b0000001b0000001b", 11674=>X"0000001b0000001b0000001b0000001b", 
11675=>X"0000001b0000001b0000001b0000001b", 11676=>X"0000001b0000001b0000001b0000001b", 11677=>X"0000001b0000001b0000001b0000001b", 11678=>X"0000001b0000001b0000001b0000001b", 11679=>X"0000001b0000001b0000001b0000001b", 
11680=>X"0000001b0000001b0000001b0000001b", 11681=>X"0000001b0000001b0000001b0000001b", 11682=>X"0000001b0000001b0000001b0000001b", 11683=>X"0000001b0000001b0000001b0000001b", 11684=>X"0000001b0000001b0000001b0000001b", 
11685=>X"0000001b0000001b0000001b0000001b", 11686=>X"0000001b0000001b0000001b0000001b", 11687=>X"0000001b0000001b0000001b0000001b", 11688=>X"0000001b0000001b0000001b0000001b", 11689=>X"0000001b0000001b0000001b0000001b", 
11690=>X"0000001b0000001b0000001b0000001b", 11691=>X"0000001b0000001b0000001b0000001b", 11692=>X"0000001b0000001b0000001b0000001b", 11693=>X"0000001b0000001b0000001b0000001b", 11694=>X"0000001b0000001b0000001b0000001b", 
11695=>X"0000001b0000001b0000001b0000001b", 11696=>X"0000001b0000001b0000001b0000001b", 11697=>X"0000001b0000001b0000001b0000001b", 11698=>X"0000001b0000001b0000001b0000001b", 11699=>X"0000001b0000001b0000001b0000001b", 
11700=>X"0000001b0000001b0000001b0000001b", 11701=>X"0000001b0000001b0000001b0000001b", 11702=>X"0000001b0000001b0000001b0000001b", 11703=>X"0000001b0000001b0000001b0000001b", 11704=>X"0000001b0000001b0000001b0000001b", 
11705=>X"0000001b0000001b0000001b0000001b", 11706=>X"0000001b0000001b0000001b0000001b", 11707=>X"0000001b0000001b0000001b0000001b", 11708=>X"0000001b0000001b0000001b0000001b", 11709=>X"0000001b0000001b0000001b0000001b", 
11710=>X"0000001b0000001b0000001b0000001b", 11711=>X"0000001b0000001b0000001b0000001b", 11712=>X"0000001b0000001b0000001b0000001b", 11713=>X"0000001b0000001b0000001b0000001b", 11714=>X"0000001b0000001b0000001b0000001b", 
11715=>X"0000001b0000001b0000001b0000001b", 11716=>X"0000001b0000001b0000001b0000001b", 11717=>X"0000001b0000001b0000001b0000001b", 11718=>X"0000001b0000001b0000001b0000001b", 11719=>X"0000001b0000001b0000001b0000001b", 
11720=>X"0000001b0000001b0000001b0000001b", 11721=>X"0000001b0000001b0000001b0000001b", 11722=>X"0000001b0000001b0000001b0000001b", 11723=>X"0000001b0000001b0000001b0000001b", 11724=>X"0000001b0000001b0000001b0000001b", 
11725=>X"0000001b0000001b0000001b0000001b", 11726=>X"0000001b0000001b0000001b0000001b", 11727=>X"0000001b0000001b0000001b0000001b", 11728=>X"0000001b0000001b0000001b0000001b", 11729=>X"0000001b0000001b0000001b0000001b", 
11730=>X"0000001b0000001b0000001b0000001b", 11731=>X"0000001b0000001b0000001b0000001b", 11732=>X"0000001b0000001b0000001b0000001b", 11733=>X"0000001b0000001b0000001b0000001b", 11734=>X"0000001b0000001b0000001b0000001b", 
11735=>X"0000001b0000001b0000001b0000001b", 11736=>X"0000001b0000001b0000001b0000001b", 11737=>X"0000001b0000001b0000001b0000001b", 11738=>X"0000001b0000001b0000001b0000001b", 11739=>X"0000001b0000001b0000001b0000001b", 
11740=>X"0000001b0000001b0000001b0000001b", 11741=>X"0000001b0000001b0000001b0000001b", 11742=>X"0000001b0000001b0000001b0000001b", 11743=>X"0000001b0000001b0000001b0000001b", 11744=>X"0000001b0000001b0000001b0000001b", 
11745=>X"0000001b0000001b0000001b0000001b", 11746=>X"0000001b0000001b0000001b0000001b", 11747=>X"0000001b0000001b0000001b0000001b", 11748=>X"0000001b0000001b0000001b0000001b", 11749=>X"0000001b0000001b0000001b0000001b", 
11750=>X"0000001b0000001b0000001b0000001b", 11751=>X"0000001b0000001b0000001b0000001b", 11752=>X"0000001b0000001b0000001b0000001b", 11753=>X"0000001b0000001b0000001b0000001b", 11754=>X"0000001b0000001b0000001b0000001b", 
11755=>X"0000001b0000001b0000001b0000001b", 11756=>X"0000001b0000001b0000001b0000001b", 11757=>X"0000001b0000001b0000001b0000001b", 11758=>X"0000001b0000001b0000001b0000001b", 11759=>X"0000001b0000001b0000001b0000001b", 
11760=>X"0000001b0000001b0000001b0000001b", 11761=>X"0000001b0000001b0000001b0000001b", 11762=>X"0000001a0000001a0000001a0000001a", 11763=>X"0000001a0000001a0000001a0000001a", 11764=>X"0000001a0000001a0000001a0000001a", 
11765=>X"0000001a0000001a0000001a0000001a", 11766=>X"0000001a0000001a0000001a0000001a", 11767=>X"0000001a0000001a0000001a0000001a", 11768=>X"0000001a0000001a0000001a0000001a", 11769=>X"0000001a0000001a0000001a0000001a", 
11770=>X"0000001a0000001a0000001a0000001a", 11771=>X"0000001a0000001a0000001a0000001a", 11772=>X"0000001a0000001a0000001a0000001a", 11773=>X"0000001a0000001a0000001a0000001a", 11774=>X"0000001a0000001a0000001a0000001a", 
11775=>X"0000001a0000001a0000001a0000001a", 11776=>X"0000001a0000001a0000001a0000001a", 11777=>X"0000001a0000001a0000001a0000001a", 11778=>X"0000001a0000001a0000001a0000001a", 11779=>X"0000001a0000001a0000001a0000001a", 
11780=>X"0000001a0000001a0000001a0000001a", 11781=>X"0000001a0000001a0000001a0000001a", 11782=>X"0000001a0000001a0000001a0000001a", 11783=>X"0000001a0000001a0000001a0000001a", 11784=>X"0000001a0000001a0000001a0000001a", 
11785=>X"0000001a0000001a0000001a0000001a", 11786=>X"0000001a0000001a0000001a0000001a", 11787=>X"0000001a0000001a0000001a0000001a", 11788=>X"0000001a0000001a0000001a0000001a", 11789=>X"0000001a0000001a0000001a0000001a", 
11790=>X"0000001a0000001a0000001a0000001a", 11791=>X"0000001a0000001a0000001a0000001a", 11792=>X"0000001a0000001a0000001a0000001a", 11793=>X"0000001a0000001a0000001a0000001a", 11794=>X"0000001a0000001a0000001a0000001a", 
11795=>X"0000001a0000001a0000001a0000001a", 11796=>X"0000001a0000001a0000001a0000001a", 11797=>X"0000001a0000001a0000001a0000001a", 11798=>X"0000001a0000001a0000001a0000001a", 11799=>X"0000001a0000001a0000001a0000001a", 
11800=>X"0000001a0000001a0000001a0000001a", 11801=>X"0000001a0000001a0000001a0000001a", 11802=>X"0000001a0000001a0000001a0000001a", 11803=>X"0000001a0000001a0000001a0000001a", 11804=>X"0000001a0000001a0000001a0000001a", 
11805=>X"0000001a0000001a0000001a0000001a", 11806=>X"0000001a0000001a0000001a0000001a", 11807=>X"0000001a0000001a0000001a0000001a", 11808=>X"0000001a0000001a0000001a0000001a", 11809=>X"0000001a0000001a0000001a0000001a", 
11810=>X"0000001a0000001a0000001a0000001a", 11811=>X"0000001a0000001a0000001a0000001a", 11812=>X"0000001a0000001a0000001a0000001a", 11813=>X"0000001a0000001a0000001a0000001a", 11814=>X"0000001a0000001a0000001a0000001a", 
11815=>X"0000001a0000001a0000001a0000001a", 11816=>X"0000001a0000001a0000001a0000001a", 11817=>X"0000001a0000001a0000001a0000001a", 11818=>X"0000001a0000001a0000001a0000001a", 11819=>X"0000001a0000001a0000001a0000001a", 
11820=>X"0000001a0000001a0000001a0000001a", 11821=>X"0000001a0000001a0000001a0000001a", 11822=>X"0000001a0000001a0000001a0000001a", 11823=>X"0000001a0000001a0000001a0000001a", 11824=>X"0000001a0000001a0000001a0000001a", 
11825=>X"0000001a0000001a0000001a0000001a", 11826=>X"0000001a0000001a0000001a0000001a", 11827=>X"0000001a0000001a0000001a0000001a", 11828=>X"0000001a0000001a0000001a0000001a", 11829=>X"0000001a0000001a0000001a0000001a", 
11830=>X"0000001a0000001a0000001a0000001a", 11831=>X"0000001a0000001a0000001a0000001a", 11832=>X"0000001a0000001a0000001a0000001a", 11833=>X"0000001a0000001a0000001a0000001a", 11834=>X"0000001a0000001a0000001a0000001a", 
11835=>X"0000001a0000001a0000001a0000001a", 11836=>X"0000001a0000001a0000001a0000001a", 11837=>X"0000001a0000001a0000001a0000001a", 11838=>X"0000001a0000001a0000001a0000001a", 11839=>X"0000001a0000001a0000001a0000001a", 
11840=>X"0000001a0000001a0000001a0000001a", 11841=>X"0000001a0000001a0000001a0000001a", 11842=>X"0000001a0000001a0000001a0000001a", 11843=>X"0000001a0000001a0000001a0000001a", 11844=>X"0000001a0000001a0000001a0000001a", 
11845=>X"0000001a0000001a0000001a0000001a", 11846=>X"0000001a0000001a0000001a0000001a", 11847=>X"0000001a0000001a0000001a0000001a", 11848=>X"0000001a0000001a0000001a0000001a", 11849=>X"0000001a0000001a0000001a0000001a", 
11850=>X"0000001a0000001a0000001a0000001a", 11851=>X"0000001a0000001a0000001a0000001a", 11852=>X"0000001a0000001a0000001a0000001a", 11853=>X"0000001a0000001a0000001a0000001a", 11854=>X"0000001a0000001a0000001a0000001a", 
11855=>X"0000001a0000001a0000001a0000001a", 11856=>X"0000001a0000001a0000001a0000001a", 11857=>X"0000001a0000001a0000001a0000001a", 11858=>X"0000001a0000001a0000001a0000001a", 11859=>X"0000001a0000001a0000001a0000001a", 
11860=>X"0000001a0000001a0000001a0000001a", 11861=>X"0000001a0000001a0000001a0000001a", 11862=>X"0000001a0000001a0000001a0000001a", 11863=>X"0000001a0000001a0000001a0000001a", 11864=>X"0000001a0000001a0000001a0000001a", 
11865=>X"0000001a0000001a0000001a0000001a", 11866=>X"0000001a0000001a0000001a0000001a", 11867=>X"0000001a0000001a0000001a0000001a", 11868=>X"0000001a0000001a0000001a0000001a", 11869=>X"0000001a0000001a0000001a0000001a", 
11870=>X"0000001a0000001a0000001a0000001a", 11871=>X"0000001a0000001a0000001a0000001a", 11872=>X"0000001a0000001a0000001a0000001a", 11873=>X"0000001a0000001a0000001a0000001a", 11874=>X"0000001a0000001a0000001a0000001a", 
11875=>X"0000001a0000001a0000001a0000001a", 11876=>X"0000001a0000001a0000001a0000001a", 11877=>X"0000001a0000001a0000001a0000001a", 11878=>X"0000001a0000001a0000001a0000001a", 11879=>X"0000001a0000001a0000001a0000001a", 
11880=>X"0000001a0000001a0000001a0000001a", 11881=>X"0000001a0000001a0000001a0000001a", 11882=>X"0000001a0000001a0000001a0000001a", 11883=>X"0000001a0000001a0000001a0000001a", 11884=>X"0000001a0000001a0000001a0000001a", 
11885=>X"0000001a0000001a0000001a0000001a", 11886=>X"0000001a0000001a0000001a0000001a", 11887=>X"0000001a0000001a0000001a0000001a", 11888=>X"0000001a0000001a0000001a0000001a", 11889=>X"0000001a0000001a0000001a0000001a", 
11890=>X"0000001a0000001a0000001a0000001a", 11891=>X"0000001a0000001a0000001a0000001a", 11892=>X"0000001a0000001a0000001a0000001a", 11893=>X"0000001a0000001a0000001a0000001a", 11894=>X"0000001a0000001a0000001a0000001a", 
11895=>X"0000001a0000001a0000001a0000001a", 11896=>X"0000001a0000001a0000001a0000001a", 11897=>X"0000001a0000001a0000001a0000001a", 11898=>X"0000001a0000001a0000001a0000001a", 11899=>X"0000001a0000001a0000001a0000001a", 
11900=>X"0000001a0000001a0000001a0000001a", 11901=>X"0000001a0000001a0000001a0000001a", 11902=>X"0000001a0000001a0000001a0000001a", 11903=>X"0000001a0000001a0000001a0000001a", 11904=>X"0000001a0000001a0000001a0000001a", 
11905=>X"0000001a0000001a0000001a0000001a", 11906=>X"0000001a0000001a0000001a0000001a", 11907=>X"0000001a0000001a0000001a0000001a", 11908=>X"0000001a0000001a0000001a0000001a", 11909=>X"0000001a0000001a0000001a0000001a", 
11910=>X"0000001a0000001a0000001a0000001a", 11911=>X"0000001a0000001a0000001a0000001a", 11912=>X"0000001a0000001a0000001a0000001a", 11913=>X"0000001a0000001a0000001a0000001a", 11914=>X"0000001a0000001a0000001a0000001a", 
11915=>X"0000001a0000001a0000001a0000001a", 11916=>X"0000001a0000001a0000001a0000001a", 11917=>X"0000001a0000001a0000001a0000001a", 11918=>X"0000001a0000001a0000001a0000001a", 11919=>X"0000001a0000001a0000001a0000001a", 
11920=>X"0000001a0000001a0000001a0000001a", 11921=>X"0000001a0000001a0000001a0000001a", 11922=>X"0000001a0000001a0000001a0000001a", 11923=>X"0000001a0000001a0000001a0000001a", 11924=>X"0000001a0000001a0000001a0000001a", 
11925=>X"0000001a0000001a0000001a0000001a", 11926=>X"0000001a0000001a0000001a0000001a", 11927=>X"0000001a0000001a0000001a0000001a", 11928=>X"0000001a0000001a0000001a0000001a", 11929=>X"0000001a0000001a0000001a0000001a", 
11930=>X"0000001a0000001a0000001a0000001a", 11931=>X"0000001a0000001a0000001a0000001a", 11932=>X"0000001a0000001a0000001a0000001a", 11933=>X"0000001a0000001a0000001a0000001a", 11934=>X"0000001a0000001a0000001a0000001a", 
11935=>X"0000001a0000001a0000001a0000001a", 11936=>X"0000001a0000001a0000001a0000001a", 11937=>X"0000001a0000001a0000001a0000001a", 11938=>X"0000001a0000001a0000001a0000001a", 11939=>X"0000001a0000001a0000001a0000001a", 
11940=>X"0000001a0000001a0000001a0000001a", 11941=>X"0000001a0000001a0000001a0000001a", 11942=>X"0000001a0000001a0000001a0000001a", 11943=>X"0000001a0000001a0000001a0000001a", 11944=>X"0000001a0000001a0000001a0000001a", 
11945=>X"0000001a0000001a0000001a0000001a", 11946=>X"0000001a0000001a0000001a0000001a", 11947=>X"0000001a0000001a0000001a0000001a", 11948=>X"0000001a0000001a0000001a0000001a", 11949=>X"0000001a0000001a0000001a0000001a", 
11950=>X"0000001a0000001a0000001a0000001a", 11951=>X"0000001a0000001a0000001a0000001a", 11952=>X"0000001a0000001a0000001a0000001a", 11953=>X"0000001a0000001a0000001a0000001a", 11954=>X"0000001a0000001a0000001a0000001a", 
11955=>X"0000001a0000001a0000001a0000001a", 11956=>X"0000001a0000001a0000001a0000001a", 11957=>X"0000001a0000001a0000001a0000001a", 11958=>X"0000001a0000001a0000001a0000001a", 11959=>X"0000001a0000001a0000001a0000001a", 
11960=>X"0000001a0000001a0000001a0000001a", 11961=>X"0000001a0000001a0000001a0000001a", 11962=>X"0000001a0000001a0000001a0000001a", 11963=>X"0000001a0000001a0000001a0000001a", 11964=>X"0000001a0000001a0000001a0000001a", 
11965=>X"0000001a0000001a0000001a0000001a", 11966=>X"0000001a0000001a0000001a0000001a", 11967=>X"0000001a0000001a0000001a0000001a", 11968=>X"0000001a0000001a0000001a0000001a", 11969=>X"0000001a0000001a0000001a0000001a", 
11970=>X"0000001a0000001a0000001a0000001a", 11971=>X"0000001a0000001a0000001a0000001a", 11972=>X"0000001a0000001a0000001a0000001a", 11973=>X"0000001a0000001a0000001a0000001a", 11974=>X"0000001a0000001a0000001a0000001a", 
11975=>X"0000001a0000001a0000001a0000001a", 11976=>X"0000001a0000001a0000001a0000001a", 11977=>X"0000001a0000001a0000001a0000001a", 11978=>X"0000001a0000001a0000001a0000001a", 11979=>X"0000001a0000001a0000001a0000001a", 
11980=>X"0000001a0000001a0000001a0000001a", 11981=>X"0000001a0000001a0000001a0000001a", 11982=>X"0000001a0000001a0000001a0000001a", 11983=>X"0000001a0000001a0000001a0000001a", 11984=>X"0000001a0000001a0000001a0000001a", 
11985=>X"0000001a0000001a0000001a0000001a", 11986=>X"0000001a0000001a0000001a0000001a", 11987=>X"0000001a0000001a0000001a0000001a", 11988=>X"0000001a0000001a0000001a0000001a", 11989=>X"0000001a0000001a0000001a0000001a", 
11990=>X"0000001a0000001a0000001a0000001a", 11991=>X"0000001a0000001a0000001a0000001a", 11992=>X"0000001a0000001a0000001a0000001a", 11993=>X"0000001a0000001a0000001a0000001a", 11994=>X"0000001a0000001a0000001a0000001a", 
11995=>X"0000001a0000001a0000001a0000001a", 11996=>X"0000001a0000001a0000001a0000001a", 11997=>X"0000001a0000001a0000001a0000001a", 11998=>X"0000001a0000001a0000001a0000001a", 11999=>X"0000001a0000001a0000001a0000001a", 
12000=>X"0000001a0000001a0000001a0000001a", 12001=>X"0000001a0000001a0000001a0000001a", 12002=>X"0000001a0000001a0000001a0000001a", 12003=>X"0000001a0000001a0000001a0000001a", 12004=>X"0000001a0000001a0000001a0000001a", 
12005=>X"0000001a0000001a0000001a0000001a", 12006=>X"0000001a0000001a0000001a0000001a", 12007=>X"0000001a0000001a0000001a0000001a", 12008=>X"0000001a0000001a0000001a0000001a", 12009=>X"0000001a0000001a0000001a0000001a", 
12010=>X"0000001a0000001a0000001a0000001a", 12011=>X"0000001a0000001a0000001a0000001a", 12012=>X"0000001a0000001a0000001a0000001a", 12013=>X"0000001a0000001a0000001a0000001a", 12014=>X"0000001a0000001a0000001a0000001a", 
12015=>X"0000001a0000001a0000001a0000001a", 12016=>X"0000001a0000001a0000001a0000001a", 12017=>X"0000001a0000001a0000001a0000001a", 12018=>X"0000001a0000001a0000001a0000001a", 12019=>X"0000001a0000001a0000001a0000001a", 
12020=>X"0000001a0000001a0000001a0000001a", 12021=>X"0000001a0000001a0000001a0000001a", 12022=>X"0000001a0000001a0000001a0000001a", 12023=>X"0000001a0000001a0000001a0000001a", 12024=>X"0000001a0000001a0000001a0000001a", 
12025=>X"0000001a0000001a0000001a0000001a", 12026=>X"0000001a0000001a0000001a0000001a", 12027=>X"0000001a0000001a0000001a0000001a", 12028=>X"0000001a0000001a0000001a0000001a", 12029=>X"0000001a0000001a0000001a0000001a", 
12030=>X"0000001a0000001a0000001a0000001a", 12031=>X"0000001a0000001a0000001a0000001a", 12032=>X"0000001a0000001a0000001a0000001a", 12033=>X"0000001a0000001a0000001a0000001a", 12034=>X"0000001a0000001a0000001a0000001a", 
12035=>X"0000001a0000001a0000001a0000001a", 12036=>X"0000001a0000001a0000001a0000001a", 12037=>X"0000001a0000001a0000001a0000001a", 12038=>X"0000001a0000001a0000001a0000001a", 12039=>X"0000001a0000001a0000001a0000001a", 
12040=>X"0000001a0000001a0000001a0000001a", 12041=>X"0000001a0000001a0000001a0000001a", 12042=>X"0000001a0000001a0000001a0000001a", 12043=>X"0000001a0000001a0000001a0000001a", 12044=>X"0000001a0000001a0000001a0000001a", 
12045=>X"0000001a0000001a0000001a0000001a", 12046=>X"0000001a0000001a0000001a0000001a", 12047=>X"0000001a0000001a0000001a0000001a", 12048=>X"0000001a0000001a0000001a0000001a", 12049=>X"0000001a0000001a0000001a0000001a", 
12050=>X"0000001a0000001a0000001a0000001a", 12051=>X"0000001a0000001a0000001a0000001a", 12052=>X"0000001a0000001a0000001a0000001a", 12053=>X"0000001a0000001a0000001a0000001a", 12054=>X"0000001a0000001a0000001a0000001a", 
12055=>X"0000001a0000001a0000001a0000001a", 12056=>X"0000001a0000001a0000001a0000001a", 12057=>X"0000001a0000001a0000001a0000001a", 12058=>X"0000001a0000001a0000001a0000001a", 12059=>X"0000001a0000001a0000001a0000001a", 
12060=>X"0000001a0000001a0000001a0000001a", 12061=>X"0000001a0000001a0000001a0000001a", 12062=>X"0000001a0000001a0000001a0000001a", 12063=>X"0000001a0000001a0000001a0000001a", 12064=>X"0000001a0000001a0000001a0000001a", 
12065=>X"0000001a0000001a0000001a0000001a", 12066=>X"0000001a0000001a0000001a0000001a", 12067=>X"0000001a0000001a0000001a0000001a", 12068=>X"0000001a0000001a0000001a0000001a", 12069=>X"0000001a0000001a0000001a0000001a", 
12070=>X"0000001a0000001a0000001a0000001a", 12071=>X"0000001a0000001a0000001a0000001a", 12072=>X"0000001a0000001a0000001a0000001a", 12073=>X"0000001a0000001a0000001a0000001a", 12074=>X"0000001a0000001a0000001a0000001a", 
12075=>X"0000001a0000001a0000001a0000001a", 12076=>X"0000001a0000001a0000001a0000001a", 12077=>X"0000001a0000001a0000001a0000001a", 12078=>X"0000001a0000001a0000001a0000001a", 12079=>X"0000001a0000001a0000001a0000001a", 
12080=>X"0000001a0000001a0000001a0000001a", 12081=>X"0000001a0000001a0000001a0000001a", 12082=>X"0000001a0000001a0000001a0000001a", 12083=>X"0000001a0000001a0000001a0000001a", 12084=>X"0000001a0000001a0000001a0000001a", 
12085=>X"0000001a0000001a0000001a0000001a", 12086=>X"0000001a0000001a0000001a0000001a", 12087=>X"0000001a0000001a0000001a0000001a", 12088=>X"0000001a0000001a0000001a0000001a", 12089=>X"0000001a0000001a0000001a0000001a", 
12090=>X"0000001a0000001a0000001a0000001a", 12091=>X"0000001a0000001a0000001a0000001a", 12092=>X"0000001a0000001a0000001a0000001a", 12093=>X"0000001a0000001a0000001a0000001a", 12094=>X"0000001a0000001a0000001a0000001a", 
12095=>X"0000001a0000001a0000001a0000001a", 12096=>X"0000001a0000001a0000001a0000001a", 12097=>X"0000001a0000001a0000001a0000001a", 12098=>X"0000001a0000001a0000001a0000001a", 12099=>X"0000001a0000001a0000001a0000001a", 
12100=>X"0000001a0000001a0000001a0000001a", 12101=>X"0000001a0000001a0000001a0000001a", 12102=>X"0000001a0000001a0000001a0000001a", 12103=>X"0000001a0000001a0000001a0000001a", 12104=>X"0000001a0000001a0000001a0000001a", 
12105=>X"0000001a0000001a0000001a0000001a", 12106=>X"0000001a0000001a0000001a0000001a", 12107=>X"0000001a0000001a0000001a0000001a", 12108=>X"0000001a0000001a0000001a0000001a", 12109=>X"0000001a0000001a0000001a0000001a", 
12110=>X"0000001a0000001a0000001a0000001a", 12111=>X"0000001a0000001a0000001a0000001a", 12112=>X"0000001a0000001a0000001a0000001a", 12113=>X"0000001a0000001a0000001a0000001a", 12114=>X"0000001a0000001a0000001a0000001a", 
12115=>X"0000001a0000001a0000001a0000001a", 12116=>X"0000001a0000001a0000001a0000001a", 12117=>X"0000001a0000001a0000001a0000001a", 12118=>X"0000001a0000001a0000001a0000001a", 12119=>X"0000001a0000001a0000001a0000001a", 
12120=>X"0000001a0000001a0000001a0000001a", 12121=>X"0000001a0000001a0000001a0000001a", 12122=>X"0000001a0000001a0000001a0000001a", 12123=>X"0000001a0000001a0000001a0000001a", 12124=>X"0000001a0000001a0000001a0000001a", 
12125=>X"0000001a0000001a0000001a0000001a", 12126=>X"0000001a0000001a0000001a0000001a", 12127=>X"0000001a0000001a0000001a0000001a", 12128=>X"0000001a0000001a0000001a0000001a", 12129=>X"0000001a0000001a0000001a0000001a", 
12130=>X"0000001a0000001a0000001a0000001a", 12131=>X"0000001a0000001a0000001a0000001a", 12132=>X"0000001a0000001a0000001a0000001a", 12133=>X"0000001a0000001a0000001a0000001a", 12134=>X"0000001a0000001a0000001a0000001a", 
12135=>X"0000001a0000001a0000001a0000001a", 12136=>X"0000001a0000001a0000001a0000001a", 12137=>X"0000001a0000001a0000001a0000001a", 12138=>X"0000001a0000001a0000001a0000001a", 12139=>X"0000001a0000001a0000001a0000001a", 
12140=>X"0000001a0000001a0000001a0000001a", 12141=>X"0000001a0000001a0000001a0000001a", 12142=>X"0000001a0000001a0000001a0000001a", 12143=>X"0000001a0000001a0000001a0000001a", 12144=>X"0000001a0000001a0000001a0000001a", 
12145=>X"0000001a0000001a0000001a0000001a", 12146=>X"0000001a0000001a0000001a0000001a", 12147=>X"0000001a0000001a0000001a0000001a", 12148=>X"0000001a0000001a0000001a0000001a", 12149=>X"0000001a0000001a0000001a0000001a", 
12150=>X"00000019000000190000001900000019", 12151=>X"00000019000000190000001900000019", 12152=>X"00000019000000190000001900000019", 12153=>X"00000019000000190000001900000019", 12154=>X"00000019000000190000001900000019", 
12155=>X"00000019000000190000001900000019", 12156=>X"00000019000000190000001900000019", 12157=>X"00000019000000190000001900000019", 12158=>X"00000019000000190000001900000019", 12159=>X"00000019000000190000001900000019", 
12160=>X"00000019000000190000001900000019", 12161=>X"00000019000000190000001900000019", 12162=>X"00000019000000190000001900000019", 12163=>X"00000019000000190000001900000019", 12164=>X"00000019000000190000001900000019", 
12165=>X"00000019000000190000001900000019", 12166=>X"00000019000000190000001900000019", 12167=>X"00000019000000190000001900000019", 12168=>X"00000019000000190000001900000019", 12169=>X"00000019000000190000001900000019", 
12170=>X"00000019000000190000001900000019", 12171=>X"00000019000000190000001900000019", 12172=>X"00000019000000190000001900000019", 12173=>X"00000019000000190000001900000019", 12174=>X"00000019000000190000001900000019", 
12175=>X"00000019000000190000001900000019", 12176=>X"00000019000000190000001900000019", 12177=>X"00000019000000190000001900000019", 12178=>X"00000019000000190000001900000019", 12179=>X"00000019000000190000001900000019", 
12180=>X"00000019000000190000001900000019", 12181=>X"00000019000000190000001900000019", 12182=>X"00000019000000190000001900000019", 12183=>X"00000019000000190000001900000019", 12184=>X"00000019000000190000001900000019", 
12185=>X"00000019000000190000001900000019", 12186=>X"00000019000000190000001900000019", 12187=>X"00000019000000190000001900000019", 12188=>X"00000019000000190000001900000019", 12189=>X"00000019000000190000001900000019", 
12190=>X"00000019000000190000001900000019", 12191=>X"00000019000000190000001900000019", 12192=>X"00000019000000190000001900000019", 12193=>X"00000019000000190000001900000019", 12194=>X"00000019000000190000001900000019", 
12195=>X"00000019000000190000001900000019", 12196=>X"00000019000000190000001900000019", 12197=>X"00000019000000190000001900000019", 12198=>X"00000019000000190000001900000019", 12199=>X"00000019000000190000001900000019", 
12200=>X"00000019000000190000001900000019", 12201=>X"00000019000000190000001900000019", 12202=>X"00000019000000190000001900000019", 12203=>X"00000019000000190000001900000019", 12204=>X"00000019000000190000001900000019", 
12205=>X"00000019000000190000001900000019", 12206=>X"00000019000000190000001900000019", 12207=>X"00000019000000190000001900000019", 12208=>X"00000019000000190000001900000019", 12209=>X"00000019000000190000001900000019", 
12210=>X"00000019000000190000001900000019", 12211=>X"00000019000000190000001900000019", 12212=>X"00000019000000190000001900000019", 12213=>X"00000019000000190000001900000019", 12214=>X"00000019000000190000001900000019", 
12215=>X"00000019000000190000001900000019", 12216=>X"00000019000000190000001900000019", 12217=>X"00000019000000190000001900000019", 12218=>X"00000019000000190000001900000019", 12219=>X"00000019000000190000001900000019", 
12220=>X"00000019000000190000001900000019", 12221=>X"00000019000000190000001900000019", 12222=>X"00000019000000190000001900000019", 12223=>X"00000019000000190000001900000019", 12224=>X"00000019000000190000001900000019", 
12225=>X"00000019000000190000001900000019", 12226=>X"00000019000000190000001900000019", 12227=>X"00000019000000190000001900000019", 12228=>X"00000019000000190000001900000019", 12229=>X"00000019000000190000001900000019", 
12230=>X"00000019000000190000001900000019", 12231=>X"00000019000000190000001900000019", 12232=>X"00000019000000190000001900000019", 12233=>X"00000019000000190000001900000019", 12234=>X"00000019000000190000001900000019", 
12235=>X"00000019000000190000001900000019", 12236=>X"00000019000000190000001900000019", 12237=>X"00000019000000190000001900000019", 12238=>X"00000019000000190000001900000019", 12239=>X"00000019000000190000001900000019", 
12240=>X"00000019000000190000001900000019", 12241=>X"00000019000000190000001900000019", 12242=>X"00000019000000190000001900000019", 12243=>X"00000019000000190000001900000019", 12244=>X"00000019000000190000001900000019", 
12245=>X"00000019000000190000001900000019", 12246=>X"00000019000000190000001900000019", 12247=>X"00000019000000190000001900000019", 12248=>X"00000019000000190000001900000019", 12249=>X"00000019000000190000001900000019", 
12250=>X"00000019000000190000001900000019", 12251=>X"00000019000000190000001900000019", 12252=>X"00000019000000190000001900000019", 12253=>X"00000019000000190000001900000019", 12254=>X"00000019000000190000001900000019", 
12255=>X"00000019000000190000001900000019", 12256=>X"00000019000000190000001900000019", 12257=>X"00000019000000190000001900000019", 12258=>X"00000019000000190000001900000019", 12259=>X"00000019000000190000001900000019", 
12260=>X"00000019000000190000001900000019", 12261=>X"00000019000000190000001900000019", 12262=>X"00000019000000190000001900000019", 12263=>X"00000019000000190000001900000019", 12264=>X"00000019000000190000001900000019", 
12265=>X"00000019000000190000001900000019", 12266=>X"00000019000000190000001900000019", 12267=>X"00000019000000190000001900000019", 12268=>X"00000019000000190000001900000019", 12269=>X"00000019000000190000001900000019", 
12270=>X"00000019000000190000001900000019", 12271=>X"00000019000000190000001900000019", 12272=>X"00000019000000190000001900000019", 12273=>X"00000019000000190000001900000019", 12274=>X"00000019000000190000001900000019", 
12275=>X"00000019000000190000001900000019", 12276=>X"00000019000000190000001900000019", 12277=>X"00000019000000190000001900000019", 12278=>X"00000019000000190000001900000019", 12279=>X"00000019000000190000001900000019", 
12280=>X"00000019000000190000001900000019", 12281=>X"00000019000000190000001900000019", 12282=>X"00000019000000190000001900000019", 12283=>X"00000019000000190000001900000019", 12284=>X"00000019000000190000001900000019", 
12285=>X"00000019000000190000001900000019", 12286=>X"00000019000000190000001900000019", 12287=>X"00000019000000190000001900000019", 12288=>X"00000019000000190000001900000019", 12289=>X"00000019000000190000001900000019", 
12290=>X"00000019000000190000001900000019", 12291=>X"00000019000000190000001900000019", 12292=>X"00000019000000190000001900000019", 12293=>X"00000019000000190000001900000019", 12294=>X"00000019000000190000001900000019", 
12295=>X"00000019000000190000001900000019", 12296=>X"00000019000000190000001900000019", 12297=>X"00000019000000190000001900000019", 12298=>X"00000019000000190000001900000019", 12299=>X"00000019000000190000001900000019", 
12300=>X"00000019000000190000001900000019", 12301=>X"00000019000000190000001900000019", 12302=>X"00000019000000190000001900000019", 12303=>X"00000019000000190000001900000019", 12304=>X"00000019000000190000001900000019", 
12305=>X"00000019000000190000001900000019", 12306=>X"00000019000000190000001900000019", 12307=>X"00000019000000190000001900000019", 12308=>X"00000019000000190000001900000019", 12309=>X"00000019000000190000001900000019", 
12310=>X"00000019000000190000001900000019", 12311=>X"00000019000000190000001900000019", 12312=>X"00000019000000190000001900000019", 12313=>X"00000019000000190000001900000019", 12314=>X"00000019000000190000001900000019", 
12315=>X"00000019000000190000001900000019", 12316=>X"00000019000000190000001900000019", 12317=>X"00000019000000190000001900000019", 12318=>X"00000019000000190000001900000019", 12319=>X"00000019000000190000001900000019", 
12320=>X"00000019000000190000001900000019", 12321=>X"00000019000000190000001900000019", 12322=>X"00000019000000190000001900000019", 12323=>X"00000019000000190000001900000019", 12324=>X"00000019000000190000001900000019", 
12325=>X"00000019000000190000001900000019", 12326=>X"00000019000000190000001900000019", 12327=>X"00000019000000190000001900000019", 12328=>X"00000019000000190000001900000019", 12329=>X"00000019000000190000001900000019", 
12330=>X"00000019000000190000001900000019", 12331=>X"00000019000000190000001900000019", 12332=>X"00000019000000190000001900000019", 12333=>X"00000019000000190000001900000019", 12334=>X"00000019000000190000001900000019", 
12335=>X"00000019000000190000001900000019", 12336=>X"00000019000000190000001900000019", 12337=>X"00000019000000190000001900000019", 12338=>X"00000019000000190000001900000019", 12339=>X"00000019000000190000001900000019", 
12340=>X"00000019000000190000001900000019", 12341=>X"00000019000000190000001900000019", 12342=>X"00000019000000190000001900000019", 12343=>X"00000019000000190000001900000019", 12344=>X"00000019000000190000001900000019", 
12345=>X"00000019000000190000001900000019", 12346=>X"00000019000000190000001900000019", 12347=>X"00000019000000190000001900000019", 12348=>X"00000019000000190000001900000019", 12349=>X"00000019000000190000001900000019", 
12350=>X"00000019000000190000001900000019", 12351=>X"00000019000000190000001900000019", 12352=>X"00000019000000190000001900000019", 12353=>X"00000019000000190000001900000019", 12354=>X"00000019000000190000001900000019", 
12355=>X"00000019000000190000001900000019", 12356=>X"00000019000000190000001900000019", 12357=>X"00000019000000190000001900000019", 12358=>X"00000019000000190000001900000019", 12359=>X"00000019000000190000001900000019", 
12360=>X"00000019000000190000001900000019", 12361=>X"00000019000000190000001900000019", 12362=>X"00000019000000190000001900000019", 12363=>X"00000019000000190000001900000019", 12364=>X"00000019000000190000001900000019", 
12365=>X"00000019000000190000001900000019", 12366=>X"00000019000000190000001900000019", 12367=>X"00000019000000190000001900000019", 12368=>X"00000019000000190000001900000019", 12369=>X"00000019000000190000001900000019", 
12370=>X"00000019000000190000001900000019", 12371=>X"00000019000000190000001900000019", 12372=>X"00000019000000190000001900000019", 12373=>X"00000019000000190000001900000019", 12374=>X"00000019000000190000001900000019", 
12375=>X"00000019000000190000001900000019", 12376=>X"00000019000000190000001900000019", 12377=>X"00000019000000190000001900000019", 12378=>X"00000019000000190000001900000019", 12379=>X"00000019000000190000001900000019", 
12380=>X"00000019000000190000001900000019", 12381=>X"00000019000000190000001900000019", 12382=>X"00000019000000190000001900000019", 12383=>X"00000019000000190000001900000019", 12384=>X"00000019000000190000001900000019", 
12385=>X"00000019000000190000001900000019", 12386=>X"00000019000000190000001900000019", 12387=>X"00000019000000190000001900000019", 12388=>X"00000019000000190000001900000019", 12389=>X"00000019000000190000001900000019", 
12390=>X"00000019000000190000001900000019", 12391=>X"00000019000000190000001900000019", 12392=>X"00000019000000190000001900000019", 12393=>X"00000019000000190000001900000019", 12394=>X"00000019000000190000001900000019", 
12395=>X"00000019000000190000001900000019", 12396=>X"00000019000000190000001900000019", 12397=>X"00000019000000190000001900000019", 12398=>X"00000019000000190000001900000019", 12399=>X"00000019000000190000001900000019", 
12400=>X"00000019000000190000001900000019", 12401=>X"00000019000000190000001900000019", 12402=>X"00000019000000190000001900000019", 12403=>X"00000019000000190000001900000019", 12404=>X"00000019000000190000001900000019", 
12405=>X"00000019000000190000001900000019", 12406=>X"00000019000000190000001900000019", 12407=>X"00000019000000190000001900000019", 12408=>X"00000019000000190000001900000019", 12409=>X"00000019000000190000001900000019", 
12410=>X"00000019000000190000001900000019", 12411=>X"00000019000000190000001900000019", 12412=>X"00000019000000190000001900000019", 12413=>X"00000019000000190000001900000019", 12414=>X"00000019000000190000001900000019", 
12415=>X"00000019000000190000001900000019", 12416=>X"00000019000000190000001900000019", 12417=>X"00000019000000190000001900000019", 12418=>X"00000019000000190000001900000019", 12419=>X"00000019000000190000001900000019", 
12420=>X"00000019000000190000001900000019", 12421=>X"00000019000000190000001900000019", 12422=>X"00000019000000190000001900000019", 12423=>X"00000019000000190000001900000019", 12424=>X"00000019000000190000001900000019", 
12425=>X"00000019000000190000001900000019", 12426=>X"00000019000000190000001900000019", 12427=>X"00000019000000190000001900000019", 12428=>X"00000019000000190000001900000019", 12429=>X"00000019000000190000001900000019", 
12430=>X"00000019000000190000001900000019", 12431=>X"00000019000000190000001900000019", 12432=>X"00000019000000190000001900000019", 12433=>X"00000019000000190000001900000019", 12434=>X"00000019000000190000001900000019", 
12435=>X"00000019000000190000001900000019", 12436=>X"00000019000000190000001900000019", 12437=>X"00000019000000190000001900000019", 12438=>X"00000019000000190000001900000019", 12439=>X"00000019000000190000001900000019", 
12440=>X"00000019000000190000001900000019", 12441=>X"00000019000000190000001900000019", 12442=>X"00000019000000190000001900000019", 12443=>X"00000019000000190000001900000019", 12444=>X"00000019000000190000001900000019", 
12445=>X"00000019000000190000001900000019", 12446=>X"00000019000000190000001900000019", 12447=>X"00000019000000190000001900000019", 12448=>X"00000019000000190000001900000019", 12449=>X"00000019000000190000001900000019", 
12450=>X"00000019000000190000001900000019", 12451=>X"00000019000000190000001900000019", 12452=>X"00000019000000190000001900000019", 12453=>X"00000019000000190000001900000019", 12454=>X"00000019000000190000001900000019", 
12455=>X"00000019000000190000001900000019", 12456=>X"00000019000000190000001900000019", 12457=>X"00000019000000190000001900000019", 12458=>X"00000019000000190000001900000019", 12459=>X"00000019000000190000001900000019", 
12460=>X"00000019000000190000001900000019", 12461=>X"00000019000000190000001900000019", 12462=>X"00000019000000190000001900000019", 12463=>X"00000019000000190000001900000019", 12464=>X"00000019000000190000001900000019", 
12465=>X"00000019000000190000001900000019", 12466=>X"00000019000000190000001900000019", 12467=>X"00000019000000190000001900000019", 12468=>X"00000019000000190000001900000019", 12469=>X"00000019000000190000001900000019", 
12470=>X"00000019000000190000001900000019", 12471=>X"00000019000000190000001900000019", 12472=>X"00000019000000190000001900000019", 12473=>X"00000019000000190000001900000019", 12474=>X"00000019000000190000001900000019", 
12475=>X"00000019000000190000001900000019", 12476=>X"00000019000000190000001900000019", 12477=>X"00000019000000190000001900000019", 12478=>X"00000019000000190000001900000019", 12479=>X"00000019000000190000001900000019", 
12480=>X"00000019000000190000001900000019", 12481=>X"00000019000000190000001900000019", 12482=>X"00000019000000190000001900000019", 12483=>X"00000019000000190000001900000019", 12484=>X"00000019000000190000001900000019", 
12485=>X"00000019000000190000001900000019", 12486=>X"00000019000000190000001900000019", 12487=>X"00000019000000190000001900000019", 12488=>X"00000019000000190000001900000019", 12489=>X"00000019000000190000001900000019", 
12490=>X"00000019000000190000001900000019", 12491=>X"00000019000000190000001900000019", 12492=>X"00000019000000190000001900000019", 12493=>X"00000019000000190000001900000019", 12494=>X"00000019000000190000001900000019", 
12495=>X"00000019000000190000001900000019", 12496=>X"00000019000000190000001900000019", 12497=>X"00000019000000190000001900000019", 12498=>X"00000019000000190000001900000019", 12499=>X"00000019000000190000001900000019", 
12500=>X"00000019000000190000001900000019", 12501=>X"00000019000000190000001900000019", 12502=>X"00000019000000190000001900000019", 12503=>X"00000019000000190000001900000019", 12504=>X"00000019000000190000001900000019", 
12505=>X"00000019000000190000001900000019", 12506=>X"00000019000000190000001900000019", 12507=>X"00000019000000190000001900000019", 12508=>X"00000019000000190000001900000019", 12509=>X"00000019000000190000001900000019", 
12510=>X"00000019000000190000001900000019", 12511=>X"00000019000000190000001900000019", 12512=>X"00000019000000190000001900000019", 12513=>X"00000019000000190000001900000019", 12514=>X"00000019000000190000001900000019", 
12515=>X"00000019000000190000001900000019", 12516=>X"00000019000000190000001900000019", 12517=>X"00000019000000190000001900000019", 12518=>X"00000019000000190000001900000019", 12519=>X"00000019000000190000001900000019", 
12520=>X"00000019000000190000001900000019", 12521=>X"00000019000000190000001900000019", 12522=>X"00000019000000190000001900000019", 12523=>X"00000019000000190000001900000019", 12524=>X"00000019000000190000001900000019", 
12525=>X"00000019000000190000001900000019", 12526=>X"00000019000000190000001900000019", 12527=>X"00000019000000190000001900000019", 12528=>X"00000019000000190000001900000019", 12529=>X"00000019000000190000001900000019", 
12530=>X"00000019000000190000001900000019", 12531=>X"00000019000000190000001900000019", 12532=>X"00000019000000190000001900000019", 12533=>X"00000019000000190000001900000019", 12534=>X"00000019000000190000001900000019", 
12535=>X"00000019000000190000001900000019", 12536=>X"00000019000000190000001900000019", 12537=>X"00000019000000190000001900000019", 12538=>X"00000019000000190000001900000019", 12539=>X"00000019000000190000001900000019", 
12540=>X"00000019000000190000001900000019", 12541=>X"00000019000000190000001900000019", 12542=>X"00000019000000190000001900000019", 12543=>X"00000019000000190000001900000019", 12544=>X"00000019000000190000001900000019", 
12545=>X"00000019000000190000001900000019", 12546=>X"00000019000000190000001900000019", 12547=>X"00000019000000190000001900000019", 12548=>X"00000019000000190000001900000019", 12549=>X"00000019000000190000001900000019", 
12550=>X"00000019000000190000001900000019", 12551=>X"00000019000000190000001900000019", 12552=>X"00000019000000190000001900000019", 12553=>X"00000019000000190000001900000019", 12554=>X"00000019000000190000001900000019", 
12555=>X"00000019000000190000001900000019", 12556=>X"00000019000000190000001900000019", 12557=>X"00000019000000190000001900000019", 12558=>X"00000019000000190000001900000019", 12559=>X"00000019000000190000001900000019", 
12560=>X"00000019000000190000001900000019", 12561=>X"00000019000000190000001900000019", 12562=>X"00000019000000190000001900000019", 12563=>X"00000019000000190000001900000019", 12564=>X"00000019000000190000001900000019", 
12565=>X"00000019000000190000001900000019", 12566=>X"00000019000000190000001900000019", 12567=>X"00000019000000190000001900000019", 12568=>X"00000019000000190000001900000019", 12569=>X"00000018000000190000001900000019", 
12570=>X"00000018000000180000001800000018", 12571=>X"00000018000000180000001800000018", 12572=>X"00000018000000180000001800000018", 12573=>X"00000018000000180000001800000018", 12574=>X"00000018000000180000001800000018", 
12575=>X"00000018000000180000001800000018", 12576=>X"00000018000000180000001800000018", 12577=>X"00000018000000180000001800000018", 12578=>X"00000018000000180000001800000018", 12579=>X"00000018000000180000001800000018", 
12580=>X"00000018000000180000001800000018", 12581=>X"00000018000000180000001800000018", 12582=>X"00000018000000180000001800000018", 12583=>X"00000018000000180000001800000018", 12584=>X"00000018000000180000001800000018", 
12585=>X"00000018000000180000001800000018", 12586=>X"00000018000000180000001800000018", 12587=>X"00000018000000180000001800000018", 12588=>X"00000018000000180000001800000018", 12589=>X"00000018000000180000001800000018", 
12590=>X"00000018000000180000001800000018", 12591=>X"00000018000000180000001800000018", 12592=>X"00000018000000180000001800000018", 12593=>X"00000018000000180000001800000018", 12594=>X"00000018000000180000001800000018", 
12595=>X"00000018000000180000001800000018", 12596=>X"00000018000000180000001800000018", 12597=>X"00000018000000180000001800000018", 12598=>X"00000018000000180000001800000018", 12599=>X"00000018000000180000001800000018", 
12600=>X"00000018000000180000001800000018", 12601=>X"00000018000000180000001800000018", 12602=>X"00000018000000180000001800000018", 12603=>X"00000018000000180000001800000018", 12604=>X"00000018000000180000001800000018", 
12605=>X"00000018000000180000001800000018", 12606=>X"00000018000000180000001800000018", 12607=>X"00000018000000180000001800000018", 12608=>X"00000018000000180000001800000018", 12609=>X"00000018000000180000001800000018", 
12610=>X"00000018000000180000001800000018", 12611=>X"00000018000000180000001800000018", 12612=>X"00000018000000180000001800000018", 12613=>X"00000018000000180000001800000018", 12614=>X"00000018000000180000001800000018", 
12615=>X"00000018000000180000001800000018", 12616=>X"00000018000000180000001800000018", 12617=>X"00000018000000180000001800000018", 12618=>X"00000018000000180000001800000018", 12619=>X"00000018000000180000001800000018", 
12620=>X"00000018000000180000001800000018", 12621=>X"00000018000000180000001800000018", 12622=>X"00000018000000180000001800000018", 12623=>X"00000018000000180000001800000018", 12624=>X"00000018000000180000001800000018", 
12625=>X"00000018000000180000001800000018", 12626=>X"00000018000000180000001800000018", 12627=>X"00000018000000180000001800000018", 12628=>X"00000018000000180000001800000018", 12629=>X"00000018000000180000001800000018", 
12630=>X"00000018000000180000001800000018", 12631=>X"00000018000000180000001800000018", 12632=>X"00000018000000180000001800000018", 12633=>X"00000018000000180000001800000018", 12634=>X"00000018000000180000001800000018", 
12635=>X"00000018000000180000001800000018", 12636=>X"00000018000000180000001800000018", 12637=>X"00000018000000180000001800000018", 12638=>X"00000018000000180000001800000018", 12639=>X"00000018000000180000001800000018", 
12640=>X"00000018000000180000001800000018", 12641=>X"00000018000000180000001800000018", 12642=>X"00000018000000180000001800000018", 12643=>X"00000018000000180000001800000018", 12644=>X"00000018000000180000001800000018", 
12645=>X"00000018000000180000001800000018", 12646=>X"00000018000000180000001800000018", 12647=>X"00000018000000180000001800000018", 12648=>X"00000018000000180000001800000018", 12649=>X"00000018000000180000001800000018", 
12650=>X"00000018000000180000001800000018", 12651=>X"00000018000000180000001800000018", 12652=>X"00000018000000180000001800000018", 12653=>X"00000018000000180000001800000018", 12654=>X"00000018000000180000001800000018", 
12655=>X"00000018000000180000001800000018", 12656=>X"00000018000000180000001800000018", 12657=>X"00000018000000180000001800000018", 12658=>X"00000018000000180000001800000018", 12659=>X"00000018000000180000001800000018", 
12660=>X"00000018000000180000001800000018", 12661=>X"00000018000000180000001800000018", 12662=>X"00000018000000180000001800000018", 12663=>X"00000018000000180000001800000018", 12664=>X"00000018000000180000001800000018", 
12665=>X"00000018000000180000001800000018", 12666=>X"00000018000000180000001800000018", 12667=>X"00000018000000180000001800000018", 12668=>X"00000018000000180000001800000018", 12669=>X"00000018000000180000001800000018", 
12670=>X"00000018000000180000001800000018", 12671=>X"00000018000000180000001800000018", 12672=>X"00000018000000180000001800000018", 12673=>X"00000018000000180000001800000018", 12674=>X"00000018000000180000001800000018", 
12675=>X"00000018000000180000001800000018", 12676=>X"00000018000000180000001800000018", 12677=>X"00000018000000180000001800000018", 12678=>X"00000018000000180000001800000018", 12679=>X"00000018000000180000001800000018", 
12680=>X"00000018000000180000001800000018", 12681=>X"00000018000000180000001800000018", 12682=>X"00000018000000180000001800000018", 12683=>X"00000018000000180000001800000018", 12684=>X"00000018000000180000001800000018", 
12685=>X"00000018000000180000001800000018", 12686=>X"00000018000000180000001800000018", 12687=>X"00000018000000180000001800000018", 12688=>X"00000018000000180000001800000018", 12689=>X"00000018000000180000001800000018", 
12690=>X"00000018000000180000001800000018", 12691=>X"00000018000000180000001800000018", 12692=>X"00000018000000180000001800000018", 12693=>X"00000018000000180000001800000018", 12694=>X"00000018000000180000001800000018", 
12695=>X"00000018000000180000001800000018", 12696=>X"00000018000000180000001800000018", 12697=>X"00000018000000180000001800000018", 12698=>X"00000018000000180000001800000018", 12699=>X"00000018000000180000001800000018", 
12700=>X"00000018000000180000001800000018", 12701=>X"00000018000000180000001800000018", 12702=>X"00000018000000180000001800000018", 12703=>X"00000018000000180000001800000018", 12704=>X"00000018000000180000001800000018", 
12705=>X"00000018000000180000001800000018", 12706=>X"00000018000000180000001800000018", 12707=>X"00000018000000180000001800000018", 12708=>X"00000018000000180000001800000018", 12709=>X"00000018000000180000001800000018", 
12710=>X"00000018000000180000001800000018", 12711=>X"00000018000000180000001800000018", 12712=>X"00000018000000180000001800000018", 12713=>X"00000018000000180000001800000018", 12714=>X"00000018000000180000001800000018", 
12715=>X"00000018000000180000001800000018", 12716=>X"00000018000000180000001800000018", 12717=>X"00000018000000180000001800000018", 12718=>X"00000018000000180000001800000018", 12719=>X"00000018000000180000001800000018", 
12720=>X"00000018000000180000001800000018", 12721=>X"00000018000000180000001800000018", 12722=>X"00000018000000180000001800000018", 12723=>X"00000018000000180000001800000018", 12724=>X"00000018000000180000001800000018", 
12725=>X"00000018000000180000001800000018", 12726=>X"00000018000000180000001800000018", 12727=>X"00000018000000180000001800000018", 12728=>X"00000018000000180000001800000018", 12729=>X"00000018000000180000001800000018", 
12730=>X"00000018000000180000001800000018", 12731=>X"00000018000000180000001800000018", 12732=>X"00000018000000180000001800000018", 12733=>X"00000018000000180000001800000018", 12734=>X"00000018000000180000001800000018", 
12735=>X"00000018000000180000001800000018", 12736=>X"00000018000000180000001800000018", 12737=>X"00000018000000180000001800000018", 12738=>X"00000018000000180000001800000018", 12739=>X"00000018000000180000001800000018", 
12740=>X"00000018000000180000001800000018", 12741=>X"00000018000000180000001800000018", 12742=>X"00000018000000180000001800000018", 12743=>X"00000018000000180000001800000018", 12744=>X"00000018000000180000001800000018", 
12745=>X"00000018000000180000001800000018", 12746=>X"00000018000000180000001800000018", 12747=>X"00000018000000180000001800000018", 12748=>X"00000018000000180000001800000018", 12749=>X"00000018000000180000001800000018", 
12750=>X"00000018000000180000001800000018", 12751=>X"00000018000000180000001800000018", 12752=>X"00000018000000180000001800000018", 12753=>X"00000018000000180000001800000018", 12754=>X"00000018000000180000001800000018", 
12755=>X"00000018000000180000001800000018", 12756=>X"00000018000000180000001800000018", 12757=>X"00000018000000180000001800000018", 12758=>X"00000018000000180000001800000018", 12759=>X"00000018000000180000001800000018", 
12760=>X"00000018000000180000001800000018", 12761=>X"00000018000000180000001800000018", 12762=>X"00000018000000180000001800000018", 12763=>X"00000018000000180000001800000018", 12764=>X"00000018000000180000001800000018", 
12765=>X"00000018000000180000001800000018", 12766=>X"00000018000000180000001800000018", 12767=>X"00000018000000180000001800000018", 12768=>X"00000018000000180000001800000018", 12769=>X"00000018000000180000001800000018", 
12770=>X"00000018000000180000001800000018", 12771=>X"00000018000000180000001800000018", 12772=>X"00000018000000180000001800000018", 12773=>X"00000018000000180000001800000018", 12774=>X"00000018000000180000001800000018", 
12775=>X"00000018000000180000001800000018", 12776=>X"00000018000000180000001800000018", 12777=>X"00000018000000180000001800000018", 12778=>X"00000018000000180000001800000018", 12779=>X"00000018000000180000001800000018", 
12780=>X"00000018000000180000001800000018", 12781=>X"00000018000000180000001800000018", 12782=>X"00000018000000180000001800000018", 12783=>X"00000018000000180000001800000018", 12784=>X"00000018000000180000001800000018", 
12785=>X"00000018000000180000001800000018", 12786=>X"00000018000000180000001800000018", 12787=>X"00000018000000180000001800000018", 12788=>X"00000018000000180000001800000018", 12789=>X"00000018000000180000001800000018", 
12790=>X"00000018000000180000001800000018", 12791=>X"00000018000000180000001800000018", 12792=>X"00000018000000180000001800000018", 12793=>X"00000018000000180000001800000018", 12794=>X"00000018000000180000001800000018", 
12795=>X"00000018000000180000001800000018", 12796=>X"00000018000000180000001800000018", 12797=>X"00000018000000180000001800000018", 12798=>X"00000018000000180000001800000018", 12799=>X"00000018000000180000001800000018", 
12800=>X"00000018000000180000001800000018", 12801=>X"00000018000000180000001800000018", 12802=>X"00000018000000180000001800000018", 12803=>X"00000018000000180000001800000018", 12804=>X"00000018000000180000001800000018", 
12805=>X"00000018000000180000001800000018", 12806=>X"00000018000000180000001800000018", 12807=>X"00000018000000180000001800000018", 12808=>X"00000018000000180000001800000018", 12809=>X"00000018000000180000001800000018", 
12810=>X"00000018000000180000001800000018", 12811=>X"00000018000000180000001800000018", 12812=>X"00000018000000180000001800000018", 12813=>X"00000018000000180000001800000018", 12814=>X"00000018000000180000001800000018", 
12815=>X"00000018000000180000001800000018", 12816=>X"00000018000000180000001800000018", 12817=>X"00000018000000180000001800000018", 12818=>X"00000018000000180000001800000018", 12819=>X"00000018000000180000001800000018", 
12820=>X"00000018000000180000001800000018", 12821=>X"00000018000000180000001800000018", 12822=>X"00000018000000180000001800000018", 12823=>X"00000018000000180000001800000018", 12824=>X"00000018000000180000001800000018", 
12825=>X"00000018000000180000001800000018", 12826=>X"00000018000000180000001800000018", 12827=>X"00000018000000180000001800000018", 12828=>X"00000018000000180000001800000018", 12829=>X"00000018000000180000001800000018", 
12830=>X"00000018000000180000001800000018", 12831=>X"00000018000000180000001800000018", 12832=>X"00000018000000180000001800000018", 12833=>X"00000018000000180000001800000018", 12834=>X"00000018000000180000001800000018", 
12835=>X"00000018000000180000001800000018", 12836=>X"00000018000000180000001800000018", 12837=>X"00000018000000180000001800000018", 12838=>X"00000018000000180000001800000018", 12839=>X"00000018000000180000001800000018", 
12840=>X"00000018000000180000001800000018", 12841=>X"00000018000000180000001800000018", 12842=>X"00000018000000180000001800000018", 12843=>X"00000018000000180000001800000018", 12844=>X"00000018000000180000001800000018", 
12845=>X"00000018000000180000001800000018", 12846=>X"00000018000000180000001800000018", 12847=>X"00000018000000180000001800000018", 12848=>X"00000018000000180000001800000018", 12849=>X"00000018000000180000001800000018", 
12850=>X"00000018000000180000001800000018", 12851=>X"00000018000000180000001800000018", 12852=>X"00000018000000180000001800000018", 12853=>X"00000018000000180000001800000018", 12854=>X"00000018000000180000001800000018", 
12855=>X"00000018000000180000001800000018", 12856=>X"00000018000000180000001800000018", 12857=>X"00000018000000180000001800000018", 12858=>X"00000018000000180000001800000018", 12859=>X"00000018000000180000001800000018", 
12860=>X"00000018000000180000001800000018", 12861=>X"00000018000000180000001800000018", 12862=>X"00000018000000180000001800000018", 12863=>X"00000018000000180000001800000018", 12864=>X"00000018000000180000001800000018", 
12865=>X"00000018000000180000001800000018", 12866=>X"00000018000000180000001800000018", 12867=>X"00000018000000180000001800000018", 12868=>X"00000018000000180000001800000018", 12869=>X"00000018000000180000001800000018", 
12870=>X"00000018000000180000001800000018", 12871=>X"00000018000000180000001800000018", 12872=>X"00000018000000180000001800000018", 12873=>X"00000018000000180000001800000018", 12874=>X"00000018000000180000001800000018", 
12875=>X"00000018000000180000001800000018", 12876=>X"00000018000000180000001800000018", 12877=>X"00000018000000180000001800000018", 12878=>X"00000018000000180000001800000018", 12879=>X"00000018000000180000001800000018", 
12880=>X"00000018000000180000001800000018", 12881=>X"00000018000000180000001800000018", 12882=>X"00000018000000180000001800000018", 12883=>X"00000018000000180000001800000018", 12884=>X"00000018000000180000001800000018", 
12885=>X"00000018000000180000001800000018", 12886=>X"00000018000000180000001800000018", 12887=>X"00000018000000180000001800000018", 12888=>X"00000018000000180000001800000018", 12889=>X"00000018000000180000001800000018", 
12890=>X"00000018000000180000001800000018", 12891=>X"00000018000000180000001800000018", 12892=>X"00000018000000180000001800000018", 12893=>X"00000018000000180000001800000018", 12894=>X"00000018000000180000001800000018", 
12895=>X"00000018000000180000001800000018", 12896=>X"00000018000000180000001800000018", 12897=>X"00000018000000180000001800000018", 12898=>X"00000018000000180000001800000018", 12899=>X"00000018000000180000001800000018", 
12900=>X"00000018000000180000001800000018", 12901=>X"00000018000000180000001800000018", 12902=>X"00000018000000180000001800000018", 12903=>X"00000018000000180000001800000018", 12904=>X"00000018000000180000001800000018", 
12905=>X"00000018000000180000001800000018", 12906=>X"00000018000000180000001800000018", 12907=>X"00000018000000180000001800000018", 12908=>X"00000018000000180000001800000018", 12909=>X"00000018000000180000001800000018", 
12910=>X"00000018000000180000001800000018", 12911=>X"00000018000000180000001800000018", 12912=>X"00000018000000180000001800000018", 12913=>X"00000018000000180000001800000018", 12914=>X"00000018000000180000001800000018", 
12915=>X"00000018000000180000001800000018", 12916=>X"00000018000000180000001800000018", 12917=>X"00000018000000180000001800000018", 12918=>X"00000018000000180000001800000018", 12919=>X"00000018000000180000001800000018", 
12920=>X"00000018000000180000001800000018", 12921=>X"00000018000000180000001800000018", 12922=>X"00000018000000180000001800000018", 12923=>X"00000018000000180000001800000018", 12924=>X"00000018000000180000001800000018", 
12925=>X"00000018000000180000001800000018", 12926=>X"00000018000000180000001800000018", 12927=>X"00000018000000180000001800000018", 12928=>X"00000018000000180000001800000018", 12929=>X"00000018000000180000001800000018", 
12930=>X"00000018000000180000001800000018", 12931=>X"00000018000000180000001800000018", 12932=>X"00000018000000180000001800000018", 12933=>X"00000018000000180000001800000018", 12934=>X"00000018000000180000001800000018", 
12935=>X"00000018000000180000001800000018", 12936=>X"00000018000000180000001800000018", 12937=>X"00000018000000180000001800000018", 12938=>X"00000018000000180000001800000018", 12939=>X"00000018000000180000001800000018", 
12940=>X"00000018000000180000001800000018", 12941=>X"00000018000000180000001800000018", 12942=>X"00000018000000180000001800000018", 12943=>X"00000018000000180000001800000018", 12944=>X"00000018000000180000001800000018", 
12945=>X"00000018000000180000001800000018", 12946=>X"00000018000000180000001800000018", 12947=>X"00000018000000180000001800000018", 12948=>X"00000018000000180000001800000018", 12949=>X"00000018000000180000001800000018", 
12950=>X"00000018000000180000001800000018", 12951=>X"00000018000000180000001800000018", 12952=>X"00000018000000180000001800000018", 12953=>X"00000018000000180000001800000018", 12954=>X"00000018000000180000001800000018", 
12955=>X"00000018000000180000001800000018", 12956=>X"00000018000000180000001800000018", 12957=>X"00000018000000180000001800000018", 12958=>X"00000018000000180000001800000018", 12959=>X"00000018000000180000001800000018", 
12960=>X"00000018000000180000001800000018", 12961=>X"00000018000000180000001800000018", 12962=>X"00000018000000180000001800000018", 12963=>X"00000018000000180000001800000018", 12964=>X"00000018000000180000001800000018", 
12965=>X"00000018000000180000001800000018", 12966=>X"00000018000000180000001800000018", 12967=>X"00000018000000180000001800000018", 12968=>X"00000018000000180000001800000018", 12969=>X"00000018000000180000001800000018", 
12970=>X"00000018000000180000001800000018", 12971=>X"00000018000000180000001800000018", 12972=>X"00000018000000180000001800000018", 12973=>X"00000018000000180000001800000018", 12974=>X"00000018000000180000001800000018", 
12975=>X"00000018000000180000001800000018", 12976=>X"00000018000000180000001800000018", 12977=>X"00000018000000180000001800000018", 12978=>X"00000018000000180000001800000018", 12979=>X"00000018000000180000001800000018", 
12980=>X"00000018000000180000001800000018", 12981=>X"00000018000000180000001800000018", 12982=>X"00000018000000180000001800000018", 12983=>X"00000018000000180000001800000018", 12984=>X"00000018000000180000001800000018", 
12985=>X"00000018000000180000001800000018", 12986=>X"00000018000000180000001800000018", 12987=>X"00000018000000180000001800000018", 12988=>X"00000018000000180000001800000018", 12989=>X"00000018000000180000001800000018", 
12990=>X"00000018000000180000001800000018", 12991=>X"00000018000000180000001800000018", 12992=>X"00000018000000180000001800000018", 12993=>X"00000018000000180000001800000018", 12994=>X"00000018000000180000001800000018", 
12995=>X"00000018000000180000001800000018", 12996=>X"00000018000000180000001800000018", 12997=>X"00000018000000180000001800000018", 12998=>X"00000018000000180000001800000018", 12999=>X"00000018000000180000001800000018", 
13000=>X"00000018000000180000001800000018", 13001=>X"00000018000000180000001800000018", 13002=>X"00000018000000180000001800000018", 13003=>X"00000018000000180000001800000018", 13004=>X"00000018000000180000001800000018", 
13005=>X"00000018000000180000001800000018", 13006=>X"00000018000000180000001800000018", 13007=>X"00000018000000180000001800000018", 13008=>X"00000018000000180000001800000018", 13009=>X"00000018000000180000001800000018", 
13010=>X"00000018000000180000001800000018", 13011=>X"00000018000000180000001800000018", 13012=>X"00000018000000180000001800000018", 13013=>X"00000018000000180000001800000018", 13014=>X"00000018000000180000001800000018", 
13015=>X"00000018000000180000001800000018", 13016=>X"00000018000000180000001800000018", 13017=>X"00000018000000180000001800000018", 13018=>X"00000018000000180000001800000018", 13019=>X"00000018000000180000001800000018", 
13020=>X"00000018000000180000001800000018", 13021=>X"00000018000000180000001800000018", 13022=>X"00000018000000180000001800000018", 13023=>X"00000018000000180000001800000018", 13024=>X"00000018000000180000001800000018", 
13025=>X"00000017000000170000001700000017", 13026=>X"00000017000000170000001700000017", 13027=>X"00000017000000170000001700000017", 13028=>X"00000017000000170000001700000017", 13029=>X"00000017000000170000001700000017", 
13030=>X"00000017000000170000001700000017", 13031=>X"00000017000000170000001700000017", 13032=>X"00000017000000170000001700000017", 13033=>X"00000017000000170000001700000017", 13034=>X"00000017000000170000001700000017", 
13035=>X"00000017000000170000001700000017", 13036=>X"00000017000000170000001700000017", 13037=>X"00000017000000170000001700000017", 13038=>X"00000017000000170000001700000017", 13039=>X"00000017000000170000001700000017", 
13040=>X"00000017000000170000001700000017", 13041=>X"00000017000000170000001700000017", 13042=>X"00000017000000170000001700000017", 13043=>X"00000017000000170000001700000017", 13044=>X"00000017000000170000001700000017", 
13045=>X"00000017000000170000001700000017", 13046=>X"00000017000000170000001700000017", 13047=>X"00000017000000170000001700000017", 13048=>X"00000017000000170000001700000017", 13049=>X"00000017000000170000001700000017", 
13050=>X"00000017000000170000001700000017", 13051=>X"00000017000000170000001700000017", 13052=>X"00000017000000170000001700000017", 13053=>X"00000017000000170000001700000017", 13054=>X"00000017000000170000001700000017", 
13055=>X"00000017000000170000001700000017", 13056=>X"00000017000000170000001700000017", 13057=>X"00000017000000170000001700000017", 13058=>X"00000017000000170000001700000017", 13059=>X"00000017000000170000001700000017", 
13060=>X"00000017000000170000001700000017", 13061=>X"00000017000000170000001700000017", 13062=>X"00000017000000170000001700000017", 13063=>X"00000017000000170000001700000017", 13064=>X"00000017000000170000001700000017", 
13065=>X"00000017000000170000001700000017", 13066=>X"00000017000000170000001700000017", 13067=>X"00000017000000170000001700000017", 13068=>X"00000017000000170000001700000017", 13069=>X"00000017000000170000001700000017", 
13070=>X"00000017000000170000001700000017", 13071=>X"00000017000000170000001700000017", 13072=>X"00000017000000170000001700000017", 13073=>X"00000017000000170000001700000017", 13074=>X"00000017000000170000001700000017", 
13075=>X"00000017000000170000001700000017", 13076=>X"00000017000000170000001700000017", 13077=>X"00000017000000170000001700000017", 13078=>X"00000017000000170000001700000017", 13079=>X"00000017000000170000001700000017", 
13080=>X"00000017000000170000001700000017", 13081=>X"00000017000000170000001700000017", 13082=>X"00000017000000170000001700000017", 13083=>X"00000017000000170000001700000017", 13084=>X"00000017000000170000001700000017", 
13085=>X"00000017000000170000001700000017", 13086=>X"00000017000000170000001700000017", 13087=>X"00000017000000170000001700000017", 13088=>X"00000017000000170000001700000017", 13089=>X"00000017000000170000001700000017", 
13090=>X"00000017000000170000001700000017", 13091=>X"00000017000000170000001700000017", 13092=>X"00000017000000170000001700000017", 13093=>X"00000017000000170000001700000017", 13094=>X"00000017000000170000001700000017", 
13095=>X"00000017000000170000001700000017", 13096=>X"00000017000000170000001700000017", 13097=>X"00000017000000170000001700000017", 13098=>X"00000017000000170000001700000017", 13099=>X"00000017000000170000001700000017", 
13100=>X"00000017000000170000001700000017", 13101=>X"00000017000000170000001700000017", 13102=>X"00000017000000170000001700000017", 13103=>X"00000017000000170000001700000017", 13104=>X"00000017000000170000001700000017", 
13105=>X"00000017000000170000001700000017", 13106=>X"00000017000000170000001700000017", 13107=>X"00000017000000170000001700000017", 13108=>X"00000017000000170000001700000017", 13109=>X"00000017000000170000001700000017", 
13110=>X"00000017000000170000001700000017", 13111=>X"00000017000000170000001700000017", 13112=>X"00000017000000170000001700000017", 13113=>X"00000017000000170000001700000017", 13114=>X"00000017000000170000001700000017", 
13115=>X"00000017000000170000001700000017", 13116=>X"00000017000000170000001700000017", 13117=>X"00000017000000170000001700000017", 13118=>X"00000017000000170000001700000017", 13119=>X"00000017000000170000001700000017", 
13120=>X"00000017000000170000001700000017", 13121=>X"00000017000000170000001700000017", 13122=>X"00000017000000170000001700000017", 13123=>X"00000017000000170000001700000017", 13124=>X"00000017000000170000001700000017", 
13125=>X"00000017000000170000001700000017", 13126=>X"00000017000000170000001700000017", 13127=>X"00000017000000170000001700000017", 13128=>X"00000017000000170000001700000017", 13129=>X"00000017000000170000001700000017", 
13130=>X"00000017000000170000001700000017", 13131=>X"00000017000000170000001700000017", 13132=>X"00000017000000170000001700000017", 13133=>X"00000017000000170000001700000017", 13134=>X"00000017000000170000001700000017", 
13135=>X"00000017000000170000001700000017", 13136=>X"00000017000000170000001700000017", 13137=>X"00000017000000170000001700000017", 13138=>X"00000017000000170000001700000017", 13139=>X"00000017000000170000001700000017", 
13140=>X"00000017000000170000001700000017", 13141=>X"00000017000000170000001700000017", 13142=>X"00000017000000170000001700000017", 13143=>X"00000017000000170000001700000017", 13144=>X"00000017000000170000001700000017", 
13145=>X"00000017000000170000001700000017", 13146=>X"00000017000000170000001700000017", 13147=>X"00000017000000170000001700000017", 13148=>X"00000017000000170000001700000017", 13149=>X"00000017000000170000001700000017", 
13150=>X"00000017000000170000001700000017", 13151=>X"00000017000000170000001700000017", 13152=>X"00000017000000170000001700000017", 13153=>X"00000017000000170000001700000017", 13154=>X"00000017000000170000001700000017", 
13155=>X"00000017000000170000001700000017", 13156=>X"00000017000000170000001700000017", 13157=>X"00000017000000170000001700000017", 13158=>X"00000017000000170000001700000017", 13159=>X"00000017000000170000001700000017", 
13160=>X"00000017000000170000001700000017", 13161=>X"00000017000000170000001700000017", 13162=>X"00000017000000170000001700000017", 13163=>X"00000017000000170000001700000017", 13164=>X"00000017000000170000001700000017", 
13165=>X"00000017000000170000001700000017", 13166=>X"00000017000000170000001700000017", 13167=>X"00000017000000170000001700000017", 13168=>X"00000017000000170000001700000017", 13169=>X"00000017000000170000001700000017", 
13170=>X"00000017000000170000001700000017", 13171=>X"00000017000000170000001700000017", 13172=>X"00000017000000170000001700000017", 13173=>X"00000017000000170000001700000017", 13174=>X"00000017000000170000001700000017", 
13175=>X"00000017000000170000001700000017", 13176=>X"00000017000000170000001700000017", 13177=>X"00000017000000170000001700000017", 13178=>X"00000017000000170000001700000017", 13179=>X"00000017000000170000001700000017", 
13180=>X"00000017000000170000001700000017", 13181=>X"00000017000000170000001700000017", 13182=>X"00000017000000170000001700000017", 13183=>X"00000017000000170000001700000017", 13184=>X"00000017000000170000001700000017", 
13185=>X"00000017000000170000001700000017", 13186=>X"00000017000000170000001700000017", 13187=>X"00000017000000170000001700000017", 13188=>X"00000017000000170000001700000017", 13189=>X"00000017000000170000001700000017", 
13190=>X"00000017000000170000001700000017", 13191=>X"00000017000000170000001700000017", 13192=>X"00000017000000170000001700000017", 13193=>X"00000017000000170000001700000017", 13194=>X"00000017000000170000001700000017", 
13195=>X"00000017000000170000001700000017", 13196=>X"00000017000000170000001700000017", 13197=>X"00000017000000170000001700000017", 13198=>X"00000017000000170000001700000017", 13199=>X"00000017000000170000001700000017", 
13200=>X"00000017000000170000001700000017", 13201=>X"00000017000000170000001700000017", 13202=>X"00000017000000170000001700000017", 13203=>X"00000017000000170000001700000017", 13204=>X"00000017000000170000001700000017", 
13205=>X"00000017000000170000001700000017", 13206=>X"00000017000000170000001700000017", 13207=>X"00000017000000170000001700000017", 13208=>X"00000017000000170000001700000017", 13209=>X"00000017000000170000001700000017", 
13210=>X"00000017000000170000001700000017", 13211=>X"00000017000000170000001700000017", 13212=>X"00000017000000170000001700000017", 13213=>X"00000017000000170000001700000017", 13214=>X"00000017000000170000001700000017", 
13215=>X"00000017000000170000001700000017", 13216=>X"00000017000000170000001700000017", 13217=>X"00000017000000170000001700000017", 13218=>X"00000017000000170000001700000017", 13219=>X"00000017000000170000001700000017", 
13220=>X"00000017000000170000001700000017", 13221=>X"00000017000000170000001700000017", 13222=>X"00000017000000170000001700000017", 13223=>X"00000017000000170000001700000017", 13224=>X"00000017000000170000001700000017", 
13225=>X"00000017000000170000001700000017", 13226=>X"00000017000000170000001700000017", 13227=>X"00000017000000170000001700000017", 13228=>X"00000017000000170000001700000017", 13229=>X"00000017000000170000001700000017", 
13230=>X"00000017000000170000001700000017", 13231=>X"00000017000000170000001700000017", 13232=>X"00000017000000170000001700000017", 13233=>X"00000017000000170000001700000017", 13234=>X"00000017000000170000001700000017", 
13235=>X"00000017000000170000001700000017", 13236=>X"00000017000000170000001700000017", 13237=>X"00000017000000170000001700000017", 13238=>X"00000017000000170000001700000017", 13239=>X"00000017000000170000001700000017", 
13240=>X"00000017000000170000001700000017", 13241=>X"00000017000000170000001700000017", 13242=>X"00000017000000170000001700000017", 13243=>X"00000017000000170000001700000017", 13244=>X"00000017000000170000001700000017", 
13245=>X"00000017000000170000001700000017", 13246=>X"00000017000000170000001700000017", 13247=>X"00000017000000170000001700000017", 13248=>X"00000017000000170000001700000017", 13249=>X"00000017000000170000001700000017", 
13250=>X"00000017000000170000001700000017", 13251=>X"00000017000000170000001700000017", 13252=>X"00000017000000170000001700000017", 13253=>X"00000017000000170000001700000017", 13254=>X"00000017000000170000001700000017", 
13255=>X"00000017000000170000001700000017", 13256=>X"00000017000000170000001700000017", 13257=>X"00000017000000170000001700000017", 13258=>X"00000017000000170000001700000017", 13259=>X"00000017000000170000001700000017", 
13260=>X"00000017000000170000001700000017", 13261=>X"00000017000000170000001700000017", 13262=>X"00000017000000170000001700000017", 13263=>X"00000017000000170000001700000017", 13264=>X"00000017000000170000001700000017", 
13265=>X"00000017000000170000001700000017", 13266=>X"00000017000000170000001700000017", 13267=>X"00000017000000170000001700000017", 13268=>X"00000017000000170000001700000017", 13269=>X"00000017000000170000001700000017", 
13270=>X"00000017000000170000001700000017", 13271=>X"00000017000000170000001700000017", 13272=>X"00000017000000170000001700000017", 13273=>X"00000017000000170000001700000017", 13274=>X"00000017000000170000001700000017", 
13275=>X"00000017000000170000001700000017", 13276=>X"00000017000000170000001700000017", 13277=>X"00000017000000170000001700000017", 13278=>X"00000017000000170000001700000017", 13279=>X"00000017000000170000001700000017", 
13280=>X"00000017000000170000001700000017", 13281=>X"00000017000000170000001700000017", 13282=>X"00000017000000170000001700000017", 13283=>X"00000017000000170000001700000017", 13284=>X"00000017000000170000001700000017", 
13285=>X"00000017000000170000001700000017", 13286=>X"00000017000000170000001700000017", 13287=>X"00000017000000170000001700000017", 13288=>X"00000017000000170000001700000017", 13289=>X"00000017000000170000001700000017", 
13290=>X"00000017000000170000001700000017", 13291=>X"00000017000000170000001700000017", 13292=>X"00000017000000170000001700000017", 13293=>X"00000017000000170000001700000017", 13294=>X"00000017000000170000001700000017", 
13295=>X"00000017000000170000001700000017", 13296=>X"00000017000000170000001700000017", 13297=>X"00000017000000170000001700000017", 13298=>X"00000017000000170000001700000017", 13299=>X"00000017000000170000001700000017", 
13300=>X"00000017000000170000001700000017", 13301=>X"00000017000000170000001700000017", 13302=>X"00000017000000170000001700000017", 13303=>X"00000017000000170000001700000017", 13304=>X"00000017000000170000001700000017", 
13305=>X"00000017000000170000001700000017", 13306=>X"00000017000000170000001700000017", 13307=>X"00000017000000170000001700000017", 13308=>X"00000017000000170000001700000017", 13309=>X"00000017000000170000001700000017", 
13310=>X"00000017000000170000001700000017", 13311=>X"00000017000000170000001700000017", 13312=>X"00000017000000170000001700000017", 13313=>X"00000017000000170000001700000017", 13314=>X"00000017000000170000001700000017", 
13315=>X"00000017000000170000001700000017", 13316=>X"00000017000000170000001700000017", 13317=>X"00000017000000170000001700000017", 13318=>X"00000017000000170000001700000017", 13319=>X"00000017000000170000001700000017", 
13320=>X"00000017000000170000001700000017", 13321=>X"00000017000000170000001700000017", 13322=>X"00000017000000170000001700000017", 13323=>X"00000017000000170000001700000017", 13324=>X"00000017000000170000001700000017", 
13325=>X"00000017000000170000001700000017", 13326=>X"00000017000000170000001700000017", 13327=>X"00000017000000170000001700000017", 13328=>X"00000017000000170000001700000017", 13329=>X"00000017000000170000001700000017", 
13330=>X"00000017000000170000001700000017", 13331=>X"00000017000000170000001700000017", 13332=>X"00000017000000170000001700000017", 13333=>X"00000017000000170000001700000017", 13334=>X"00000017000000170000001700000017", 
13335=>X"00000017000000170000001700000017", 13336=>X"00000017000000170000001700000017", 13337=>X"00000017000000170000001700000017", 13338=>X"00000017000000170000001700000017", 13339=>X"00000017000000170000001700000017", 
13340=>X"00000017000000170000001700000017", 13341=>X"00000017000000170000001700000017", 13342=>X"00000017000000170000001700000017", 13343=>X"00000017000000170000001700000017", 13344=>X"00000017000000170000001700000017", 
13345=>X"00000017000000170000001700000017", 13346=>X"00000017000000170000001700000017", 13347=>X"00000017000000170000001700000017", 13348=>X"00000017000000170000001700000017", 13349=>X"00000017000000170000001700000017", 
13350=>X"00000017000000170000001700000017", 13351=>X"00000017000000170000001700000017", 13352=>X"00000017000000170000001700000017", 13353=>X"00000017000000170000001700000017", 13354=>X"00000017000000170000001700000017", 
13355=>X"00000017000000170000001700000017", 13356=>X"00000017000000170000001700000017", 13357=>X"00000017000000170000001700000017", 13358=>X"00000017000000170000001700000017", 13359=>X"00000017000000170000001700000017", 
13360=>X"00000017000000170000001700000017", 13361=>X"00000017000000170000001700000017", 13362=>X"00000017000000170000001700000017", 13363=>X"00000017000000170000001700000017", 13364=>X"00000017000000170000001700000017", 
13365=>X"00000017000000170000001700000017", 13366=>X"00000017000000170000001700000017", 13367=>X"00000017000000170000001700000017", 13368=>X"00000017000000170000001700000017", 13369=>X"00000017000000170000001700000017", 
13370=>X"00000017000000170000001700000017", 13371=>X"00000017000000170000001700000017", 13372=>X"00000017000000170000001700000017", 13373=>X"00000017000000170000001700000017", 13374=>X"00000017000000170000001700000017", 
13375=>X"00000017000000170000001700000017", 13376=>X"00000017000000170000001700000017", 13377=>X"00000017000000170000001700000017", 13378=>X"00000017000000170000001700000017", 13379=>X"00000017000000170000001700000017", 
13380=>X"00000017000000170000001700000017", 13381=>X"00000017000000170000001700000017", 13382=>X"00000017000000170000001700000017", 13383=>X"00000017000000170000001700000017", 13384=>X"00000017000000170000001700000017", 
13385=>X"00000017000000170000001700000017", 13386=>X"00000017000000170000001700000017", 13387=>X"00000017000000170000001700000017", 13388=>X"00000017000000170000001700000017", 13389=>X"00000017000000170000001700000017", 
13390=>X"00000017000000170000001700000017", 13391=>X"00000017000000170000001700000017", 13392=>X"00000017000000170000001700000017", 13393=>X"00000017000000170000001700000017", 13394=>X"00000017000000170000001700000017", 
13395=>X"00000017000000170000001700000017", 13396=>X"00000017000000170000001700000017", 13397=>X"00000017000000170000001700000017", 13398=>X"00000017000000170000001700000017", 13399=>X"00000017000000170000001700000017", 
13400=>X"00000017000000170000001700000017", 13401=>X"00000017000000170000001700000017", 13402=>X"00000017000000170000001700000017", 13403=>X"00000017000000170000001700000017", 13404=>X"00000017000000170000001700000017", 
13405=>X"00000017000000170000001700000017", 13406=>X"00000017000000170000001700000017", 13407=>X"00000017000000170000001700000017", 13408=>X"00000017000000170000001700000017", 13409=>X"00000017000000170000001700000017", 
13410=>X"00000017000000170000001700000017", 13411=>X"00000017000000170000001700000017", 13412=>X"00000017000000170000001700000017", 13413=>X"00000017000000170000001700000017", 13414=>X"00000017000000170000001700000017", 
13415=>X"00000017000000170000001700000017", 13416=>X"00000017000000170000001700000017", 13417=>X"00000017000000170000001700000017", 13418=>X"00000017000000170000001700000017", 13419=>X"00000017000000170000001700000017", 
13420=>X"00000017000000170000001700000017", 13421=>X"00000017000000170000001700000017", 13422=>X"00000017000000170000001700000017", 13423=>X"00000017000000170000001700000017", 13424=>X"00000017000000170000001700000017", 
13425=>X"00000017000000170000001700000017", 13426=>X"00000017000000170000001700000017", 13427=>X"00000017000000170000001700000017", 13428=>X"00000017000000170000001700000017", 13429=>X"00000017000000170000001700000017", 
13430=>X"00000017000000170000001700000017", 13431=>X"00000017000000170000001700000017", 13432=>X"00000017000000170000001700000017", 13433=>X"00000017000000170000001700000017", 13434=>X"00000017000000170000001700000017", 
13435=>X"00000017000000170000001700000017", 13436=>X"00000017000000170000001700000017", 13437=>X"00000017000000170000001700000017", 13438=>X"00000017000000170000001700000017", 13439=>X"00000017000000170000001700000017", 
13440=>X"00000017000000170000001700000017", 13441=>X"00000017000000170000001700000017", 13442=>X"00000017000000170000001700000017", 13443=>X"00000017000000170000001700000017", 13444=>X"00000017000000170000001700000017", 
13445=>X"00000017000000170000001700000017", 13446=>X"00000017000000170000001700000017", 13447=>X"00000017000000170000001700000017", 13448=>X"00000017000000170000001700000017", 13449=>X"00000017000000170000001700000017", 
13450=>X"00000017000000170000001700000017", 13451=>X"00000017000000170000001700000017", 13452=>X"00000017000000170000001700000017", 13453=>X"00000017000000170000001700000017", 13454=>X"00000017000000170000001700000017", 
13455=>X"00000017000000170000001700000017", 13456=>X"00000017000000170000001700000017", 13457=>X"00000017000000170000001700000017", 13458=>X"00000017000000170000001700000017", 13459=>X"00000017000000170000001700000017", 
13460=>X"00000017000000170000001700000017", 13461=>X"00000017000000170000001700000017", 13462=>X"00000017000000170000001700000017", 13463=>X"00000017000000170000001700000017", 13464=>X"00000017000000170000001700000017", 
13465=>X"00000017000000170000001700000017", 13466=>X"00000017000000170000001700000017", 13467=>X"00000017000000170000001700000017", 13468=>X"00000017000000170000001700000017", 13469=>X"00000017000000170000001700000017", 
13470=>X"00000017000000170000001700000017", 13471=>X"00000017000000170000001700000017", 13472=>X"00000017000000170000001700000017", 13473=>X"00000017000000170000001700000017", 13474=>X"00000017000000170000001700000017", 
13475=>X"00000017000000170000001700000017", 13476=>X"00000017000000170000001700000017", 13477=>X"00000017000000170000001700000017", 13478=>X"00000017000000170000001700000017", 13479=>X"00000017000000170000001700000017", 
13480=>X"00000017000000170000001700000017", 13481=>X"00000017000000170000001700000017", 13482=>X"00000017000000170000001700000017", 13483=>X"00000017000000170000001700000017", 13484=>X"00000017000000170000001700000017", 
13485=>X"00000017000000170000001700000017", 13486=>X"00000017000000170000001700000017", 13487=>X"00000017000000170000001700000017", 13488=>X"00000017000000170000001700000017", 13489=>X"00000017000000170000001700000017", 
13490=>X"00000017000000170000001700000017", 13491=>X"00000017000000170000001700000017", 13492=>X"00000017000000170000001700000017", 13493=>X"00000017000000170000001700000017", 13494=>X"00000017000000170000001700000017", 
13495=>X"00000017000000170000001700000017", 13496=>X"00000017000000170000001700000017", 13497=>X"00000017000000170000001700000017", 13498=>X"00000017000000170000001700000017", 13499=>X"00000017000000170000001700000017", 
13500=>X"00000017000000170000001700000017", 13501=>X"00000017000000170000001700000017", 13502=>X"00000017000000170000001700000017", 13503=>X"00000017000000170000001700000017", 13504=>X"00000017000000170000001700000017", 
13505=>X"00000017000000170000001700000017", 13506=>X"00000017000000170000001700000017", 13507=>X"00000017000000170000001700000017", 13508=>X"00000017000000170000001700000017", 13509=>X"00000017000000170000001700000017", 
13510=>X"00000017000000170000001700000017", 13511=>X"00000017000000170000001700000017", 13512=>X"00000017000000170000001700000017", 13513=>X"00000017000000170000001700000017", 13514=>X"00000017000000170000001700000017", 
13515=>X"00000017000000170000001700000017", 13516=>X"00000017000000170000001700000017", 13517=>X"00000017000000170000001700000017", 13518=>X"00000017000000170000001700000017", 13519=>X"00000017000000170000001700000017", 
13520=>X"00000016000000170000001700000017", 13521=>X"00000016000000160000001600000016", 13522=>X"00000016000000160000001600000016", 13523=>X"00000016000000160000001600000016", 13524=>X"00000016000000160000001600000016", 
13525=>X"00000016000000160000001600000016", 13526=>X"00000016000000160000001600000016", 13527=>X"00000016000000160000001600000016", 13528=>X"00000016000000160000001600000016", 13529=>X"00000016000000160000001600000016", 
13530=>X"00000016000000160000001600000016", 13531=>X"00000016000000160000001600000016", 13532=>X"00000016000000160000001600000016", 13533=>X"00000016000000160000001600000016", 13534=>X"00000016000000160000001600000016", 
13535=>X"00000016000000160000001600000016", 13536=>X"00000016000000160000001600000016", 13537=>X"00000016000000160000001600000016", 13538=>X"00000016000000160000001600000016", 13539=>X"00000016000000160000001600000016", 
13540=>X"00000016000000160000001600000016", 13541=>X"00000016000000160000001600000016", 13542=>X"00000016000000160000001600000016", 13543=>X"00000016000000160000001600000016", 13544=>X"00000016000000160000001600000016", 
13545=>X"00000016000000160000001600000016", 13546=>X"00000016000000160000001600000016", 13547=>X"00000016000000160000001600000016", 13548=>X"00000016000000160000001600000016", 13549=>X"00000016000000160000001600000016", 
13550=>X"00000016000000160000001600000016", 13551=>X"00000016000000160000001600000016", 13552=>X"00000016000000160000001600000016", 13553=>X"00000016000000160000001600000016", 13554=>X"00000016000000160000001600000016", 
13555=>X"00000016000000160000001600000016", 13556=>X"00000016000000160000001600000016", 13557=>X"00000016000000160000001600000016", 13558=>X"00000016000000160000001600000016", 13559=>X"00000016000000160000001600000016", 
13560=>X"00000016000000160000001600000016", 13561=>X"00000016000000160000001600000016", 13562=>X"00000016000000160000001600000016", 13563=>X"00000016000000160000001600000016", 13564=>X"00000016000000160000001600000016", 
13565=>X"00000016000000160000001600000016", 13566=>X"00000016000000160000001600000016", 13567=>X"00000016000000160000001600000016", 13568=>X"00000016000000160000001600000016", 13569=>X"00000016000000160000001600000016", 
13570=>X"00000016000000160000001600000016", 13571=>X"00000016000000160000001600000016", 13572=>X"00000016000000160000001600000016", 13573=>X"00000016000000160000001600000016", 13574=>X"00000016000000160000001600000016", 
13575=>X"00000016000000160000001600000016", 13576=>X"00000016000000160000001600000016", 13577=>X"00000016000000160000001600000016", 13578=>X"00000016000000160000001600000016", 13579=>X"00000016000000160000001600000016", 
13580=>X"00000016000000160000001600000016", 13581=>X"00000016000000160000001600000016", 13582=>X"00000016000000160000001600000016", 13583=>X"00000016000000160000001600000016", 13584=>X"00000016000000160000001600000016", 
13585=>X"00000016000000160000001600000016", 13586=>X"00000016000000160000001600000016", 13587=>X"00000016000000160000001600000016", 13588=>X"00000016000000160000001600000016", 13589=>X"00000016000000160000001600000016", 
13590=>X"00000016000000160000001600000016", 13591=>X"00000016000000160000001600000016", 13592=>X"00000016000000160000001600000016", 13593=>X"00000016000000160000001600000016", 13594=>X"00000016000000160000001600000016", 
13595=>X"00000016000000160000001600000016", 13596=>X"00000016000000160000001600000016", 13597=>X"00000016000000160000001600000016", 13598=>X"00000016000000160000001600000016", 13599=>X"00000016000000160000001600000016", 
13600=>X"00000016000000160000001600000016", 13601=>X"00000016000000160000001600000016", 13602=>X"00000016000000160000001600000016", 13603=>X"00000016000000160000001600000016", 13604=>X"00000016000000160000001600000016", 
13605=>X"00000016000000160000001600000016", 13606=>X"00000016000000160000001600000016", 13607=>X"00000016000000160000001600000016", 13608=>X"00000016000000160000001600000016", 13609=>X"00000016000000160000001600000016", 
13610=>X"00000016000000160000001600000016", 13611=>X"00000016000000160000001600000016", 13612=>X"00000016000000160000001600000016", 13613=>X"00000016000000160000001600000016", 13614=>X"00000016000000160000001600000016", 
13615=>X"00000016000000160000001600000016", 13616=>X"00000016000000160000001600000016", 13617=>X"00000016000000160000001600000016", 13618=>X"00000016000000160000001600000016", 13619=>X"00000016000000160000001600000016", 
13620=>X"00000016000000160000001600000016", 13621=>X"00000016000000160000001600000016", 13622=>X"00000016000000160000001600000016", 13623=>X"00000016000000160000001600000016", 13624=>X"00000016000000160000001600000016", 
13625=>X"00000016000000160000001600000016", 13626=>X"00000016000000160000001600000016", 13627=>X"00000016000000160000001600000016", 13628=>X"00000016000000160000001600000016", 13629=>X"00000016000000160000001600000016", 
13630=>X"00000016000000160000001600000016", 13631=>X"00000016000000160000001600000016", 13632=>X"00000016000000160000001600000016", 13633=>X"00000016000000160000001600000016", 13634=>X"00000016000000160000001600000016", 
13635=>X"00000016000000160000001600000016", 13636=>X"00000016000000160000001600000016", 13637=>X"00000016000000160000001600000016", 13638=>X"00000016000000160000001600000016", 13639=>X"00000016000000160000001600000016", 
13640=>X"00000016000000160000001600000016", 13641=>X"00000016000000160000001600000016", 13642=>X"00000016000000160000001600000016", 13643=>X"00000016000000160000001600000016", 13644=>X"00000016000000160000001600000016", 
13645=>X"00000016000000160000001600000016", 13646=>X"00000016000000160000001600000016", 13647=>X"00000016000000160000001600000016", 13648=>X"00000016000000160000001600000016", 13649=>X"00000016000000160000001600000016", 
13650=>X"00000016000000160000001600000016", 13651=>X"00000016000000160000001600000016", 13652=>X"00000016000000160000001600000016", 13653=>X"00000016000000160000001600000016", 13654=>X"00000016000000160000001600000016", 
13655=>X"00000016000000160000001600000016", 13656=>X"00000016000000160000001600000016", 13657=>X"00000016000000160000001600000016", 13658=>X"00000016000000160000001600000016", 13659=>X"00000016000000160000001600000016", 
13660=>X"00000016000000160000001600000016", 13661=>X"00000016000000160000001600000016", 13662=>X"00000016000000160000001600000016", 13663=>X"00000016000000160000001600000016", 13664=>X"00000016000000160000001600000016", 
13665=>X"00000016000000160000001600000016", 13666=>X"00000016000000160000001600000016", 13667=>X"00000016000000160000001600000016", 13668=>X"00000016000000160000001600000016", 13669=>X"00000016000000160000001600000016", 
13670=>X"00000016000000160000001600000016", 13671=>X"00000016000000160000001600000016", 13672=>X"00000016000000160000001600000016", 13673=>X"00000016000000160000001600000016", 13674=>X"00000016000000160000001600000016", 
13675=>X"00000016000000160000001600000016", 13676=>X"00000016000000160000001600000016", 13677=>X"00000016000000160000001600000016", 13678=>X"00000016000000160000001600000016", 13679=>X"00000016000000160000001600000016", 
13680=>X"00000016000000160000001600000016", 13681=>X"00000016000000160000001600000016", 13682=>X"00000016000000160000001600000016", 13683=>X"00000016000000160000001600000016", 13684=>X"00000016000000160000001600000016", 
13685=>X"00000016000000160000001600000016", 13686=>X"00000016000000160000001600000016", 13687=>X"00000016000000160000001600000016", 13688=>X"00000016000000160000001600000016", 13689=>X"00000016000000160000001600000016", 
13690=>X"00000016000000160000001600000016", 13691=>X"00000016000000160000001600000016", 13692=>X"00000016000000160000001600000016", 13693=>X"00000016000000160000001600000016", 13694=>X"00000016000000160000001600000016", 
13695=>X"00000016000000160000001600000016", 13696=>X"00000016000000160000001600000016", 13697=>X"00000016000000160000001600000016", 13698=>X"00000016000000160000001600000016", 13699=>X"00000016000000160000001600000016", 
13700=>X"00000016000000160000001600000016", 13701=>X"00000016000000160000001600000016", 13702=>X"00000016000000160000001600000016", 13703=>X"00000016000000160000001600000016", 13704=>X"00000016000000160000001600000016", 
13705=>X"00000016000000160000001600000016", 13706=>X"00000016000000160000001600000016", 13707=>X"00000016000000160000001600000016", 13708=>X"00000016000000160000001600000016", 13709=>X"00000016000000160000001600000016", 
13710=>X"00000016000000160000001600000016", 13711=>X"00000016000000160000001600000016", 13712=>X"00000016000000160000001600000016", 13713=>X"00000016000000160000001600000016", 13714=>X"00000016000000160000001600000016", 
13715=>X"00000016000000160000001600000016", 13716=>X"00000016000000160000001600000016", 13717=>X"00000016000000160000001600000016", 13718=>X"00000016000000160000001600000016", 13719=>X"00000016000000160000001600000016", 
13720=>X"00000016000000160000001600000016", 13721=>X"00000016000000160000001600000016", 13722=>X"00000016000000160000001600000016", 13723=>X"00000016000000160000001600000016", 13724=>X"00000016000000160000001600000016", 
13725=>X"00000016000000160000001600000016", 13726=>X"00000016000000160000001600000016", 13727=>X"00000016000000160000001600000016", 13728=>X"00000016000000160000001600000016", 13729=>X"00000016000000160000001600000016", 
13730=>X"00000016000000160000001600000016", 13731=>X"00000016000000160000001600000016", 13732=>X"00000016000000160000001600000016", 13733=>X"00000016000000160000001600000016", 13734=>X"00000016000000160000001600000016", 
13735=>X"00000016000000160000001600000016", 13736=>X"00000016000000160000001600000016", 13737=>X"00000016000000160000001600000016", 13738=>X"00000016000000160000001600000016", 13739=>X"00000016000000160000001600000016", 
13740=>X"00000016000000160000001600000016", 13741=>X"00000016000000160000001600000016", 13742=>X"00000016000000160000001600000016", 13743=>X"00000016000000160000001600000016", 13744=>X"00000016000000160000001600000016", 
13745=>X"00000016000000160000001600000016", 13746=>X"00000016000000160000001600000016", 13747=>X"00000016000000160000001600000016", 13748=>X"00000016000000160000001600000016", 13749=>X"00000016000000160000001600000016", 
13750=>X"00000016000000160000001600000016", 13751=>X"00000016000000160000001600000016", 13752=>X"00000016000000160000001600000016", 13753=>X"00000016000000160000001600000016", 13754=>X"00000016000000160000001600000016", 
13755=>X"00000016000000160000001600000016", 13756=>X"00000016000000160000001600000016", 13757=>X"00000016000000160000001600000016", 13758=>X"00000016000000160000001600000016", 13759=>X"00000016000000160000001600000016", 
13760=>X"00000016000000160000001600000016", 13761=>X"00000016000000160000001600000016", 13762=>X"00000016000000160000001600000016", 13763=>X"00000016000000160000001600000016", 13764=>X"00000016000000160000001600000016", 
13765=>X"00000016000000160000001600000016", 13766=>X"00000016000000160000001600000016", 13767=>X"00000016000000160000001600000016", 13768=>X"00000016000000160000001600000016", 13769=>X"00000016000000160000001600000016", 
13770=>X"00000016000000160000001600000016", 13771=>X"00000016000000160000001600000016", 13772=>X"00000016000000160000001600000016", 13773=>X"00000016000000160000001600000016", 13774=>X"00000016000000160000001600000016", 
13775=>X"00000016000000160000001600000016", 13776=>X"00000016000000160000001600000016", 13777=>X"00000016000000160000001600000016", 13778=>X"00000016000000160000001600000016", 13779=>X"00000016000000160000001600000016", 
13780=>X"00000016000000160000001600000016", 13781=>X"00000016000000160000001600000016", 13782=>X"00000016000000160000001600000016", 13783=>X"00000016000000160000001600000016", 13784=>X"00000016000000160000001600000016", 
13785=>X"00000016000000160000001600000016", 13786=>X"00000016000000160000001600000016", 13787=>X"00000016000000160000001600000016", 13788=>X"00000016000000160000001600000016", 13789=>X"00000016000000160000001600000016", 
13790=>X"00000016000000160000001600000016", 13791=>X"00000016000000160000001600000016", 13792=>X"00000016000000160000001600000016", 13793=>X"00000016000000160000001600000016", 13794=>X"00000016000000160000001600000016", 
13795=>X"00000016000000160000001600000016", 13796=>X"00000016000000160000001600000016", 13797=>X"00000016000000160000001600000016", 13798=>X"00000016000000160000001600000016", 13799=>X"00000016000000160000001600000016", 
13800=>X"00000016000000160000001600000016", 13801=>X"00000016000000160000001600000016", 13802=>X"00000016000000160000001600000016", 13803=>X"00000016000000160000001600000016", 13804=>X"00000016000000160000001600000016", 
13805=>X"00000016000000160000001600000016", 13806=>X"00000016000000160000001600000016", 13807=>X"00000016000000160000001600000016", 13808=>X"00000016000000160000001600000016", 13809=>X"00000016000000160000001600000016", 
13810=>X"00000016000000160000001600000016", 13811=>X"00000016000000160000001600000016", 13812=>X"00000016000000160000001600000016", 13813=>X"00000016000000160000001600000016", 13814=>X"00000016000000160000001600000016", 
13815=>X"00000016000000160000001600000016", 13816=>X"00000016000000160000001600000016", 13817=>X"00000016000000160000001600000016", 13818=>X"00000016000000160000001600000016", 13819=>X"00000016000000160000001600000016", 
13820=>X"00000016000000160000001600000016", 13821=>X"00000016000000160000001600000016", 13822=>X"00000016000000160000001600000016", 13823=>X"00000016000000160000001600000016", 13824=>X"00000016000000160000001600000016", 
13825=>X"00000016000000160000001600000016", 13826=>X"00000016000000160000001600000016", 13827=>X"00000016000000160000001600000016", 13828=>X"00000016000000160000001600000016", 13829=>X"00000016000000160000001600000016", 
13830=>X"00000016000000160000001600000016", 13831=>X"00000016000000160000001600000016", 13832=>X"00000016000000160000001600000016", 13833=>X"00000016000000160000001600000016", 13834=>X"00000016000000160000001600000016", 
13835=>X"00000016000000160000001600000016", 13836=>X"00000016000000160000001600000016", 13837=>X"00000016000000160000001600000016", 13838=>X"00000016000000160000001600000016", 13839=>X"00000016000000160000001600000016", 
13840=>X"00000016000000160000001600000016", 13841=>X"00000016000000160000001600000016", 13842=>X"00000016000000160000001600000016", 13843=>X"00000016000000160000001600000016", 13844=>X"00000016000000160000001600000016", 
13845=>X"00000016000000160000001600000016", 13846=>X"00000016000000160000001600000016", 13847=>X"00000016000000160000001600000016", 13848=>X"00000016000000160000001600000016", 13849=>X"00000016000000160000001600000016", 
13850=>X"00000016000000160000001600000016", 13851=>X"00000016000000160000001600000016", 13852=>X"00000016000000160000001600000016", 13853=>X"00000016000000160000001600000016", 13854=>X"00000016000000160000001600000016", 
13855=>X"00000016000000160000001600000016", 13856=>X"00000016000000160000001600000016", 13857=>X"00000016000000160000001600000016", 13858=>X"00000016000000160000001600000016", 13859=>X"00000016000000160000001600000016", 
13860=>X"00000016000000160000001600000016", 13861=>X"00000016000000160000001600000016", 13862=>X"00000016000000160000001600000016", 13863=>X"00000016000000160000001600000016", 13864=>X"00000016000000160000001600000016", 
13865=>X"00000016000000160000001600000016", 13866=>X"00000016000000160000001600000016", 13867=>X"00000016000000160000001600000016", 13868=>X"00000016000000160000001600000016", 13869=>X"00000016000000160000001600000016", 
13870=>X"00000016000000160000001600000016", 13871=>X"00000016000000160000001600000016", 13872=>X"00000016000000160000001600000016", 13873=>X"00000016000000160000001600000016", 13874=>X"00000016000000160000001600000016", 
13875=>X"00000016000000160000001600000016", 13876=>X"00000016000000160000001600000016", 13877=>X"00000016000000160000001600000016", 13878=>X"00000016000000160000001600000016", 13879=>X"00000016000000160000001600000016", 
13880=>X"00000016000000160000001600000016", 13881=>X"00000016000000160000001600000016", 13882=>X"00000016000000160000001600000016", 13883=>X"00000016000000160000001600000016", 13884=>X"00000016000000160000001600000016", 
13885=>X"00000016000000160000001600000016", 13886=>X"00000016000000160000001600000016", 13887=>X"00000016000000160000001600000016", 13888=>X"00000016000000160000001600000016", 13889=>X"00000016000000160000001600000016", 
13890=>X"00000016000000160000001600000016", 13891=>X"00000016000000160000001600000016", 13892=>X"00000016000000160000001600000016", 13893=>X"00000016000000160000001600000016", 13894=>X"00000016000000160000001600000016", 
13895=>X"00000016000000160000001600000016", 13896=>X"00000016000000160000001600000016", 13897=>X"00000016000000160000001600000016", 13898=>X"00000016000000160000001600000016", 13899=>X"00000016000000160000001600000016", 
13900=>X"00000016000000160000001600000016", 13901=>X"00000016000000160000001600000016", 13902=>X"00000016000000160000001600000016", 13903=>X"00000016000000160000001600000016", 13904=>X"00000016000000160000001600000016", 
13905=>X"00000016000000160000001600000016", 13906=>X"00000016000000160000001600000016", 13907=>X"00000016000000160000001600000016", 13908=>X"00000016000000160000001600000016", 13909=>X"00000016000000160000001600000016", 
13910=>X"00000016000000160000001600000016", 13911=>X"00000016000000160000001600000016", 13912=>X"00000016000000160000001600000016", 13913=>X"00000016000000160000001600000016", 13914=>X"00000016000000160000001600000016", 
13915=>X"00000016000000160000001600000016", 13916=>X"00000016000000160000001600000016", 13917=>X"00000016000000160000001600000016", 13918=>X"00000016000000160000001600000016", 13919=>X"00000016000000160000001600000016", 
13920=>X"00000016000000160000001600000016", 13921=>X"00000016000000160000001600000016", 13922=>X"00000016000000160000001600000016", 13923=>X"00000016000000160000001600000016", 13924=>X"00000016000000160000001600000016", 
13925=>X"00000016000000160000001600000016", 13926=>X"00000016000000160000001600000016", 13927=>X"00000016000000160000001600000016", 13928=>X"00000016000000160000001600000016", 13929=>X"00000016000000160000001600000016", 
13930=>X"00000016000000160000001600000016", 13931=>X"00000016000000160000001600000016", 13932=>X"00000016000000160000001600000016", 13933=>X"00000016000000160000001600000016", 13934=>X"00000016000000160000001600000016", 
13935=>X"00000016000000160000001600000016", 13936=>X"00000016000000160000001600000016", 13937=>X"00000016000000160000001600000016", 13938=>X"00000016000000160000001600000016", 13939=>X"00000016000000160000001600000016", 
13940=>X"00000016000000160000001600000016", 13941=>X"00000016000000160000001600000016", 13942=>X"00000016000000160000001600000016", 13943=>X"00000016000000160000001600000016", 13944=>X"00000016000000160000001600000016", 
13945=>X"00000016000000160000001600000016", 13946=>X"00000016000000160000001600000016", 13947=>X"00000016000000160000001600000016", 13948=>X"00000016000000160000001600000016", 13949=>X"00000016000000160000001600000016", 
13950=>X"00000016000000160000001600000016", 13951=>X"00000016000000160000001600000016", 13952=>X"00000016000000160000001600000016", 13953=>X"00000016000000160000001600000016", 13954=>X"00000016000000160000001600000016", 
13955=>X"00000016000000160000001600000016", 13956=>X"00000016000000160000001600000016", 13957=>X"00000016000000160000001600000016", 13958=>X"00000016000000160000001600000016", 13959=>X"00000016000000160000001600000016", 
13960=>X"00000016000000160000001600000016", 13961=>X"00000016000000160000001600000016", 13962=>X"00000016000000160000001600000016", 13963=>X"00000016000000160000001600000016", 13964=>X"00000016000000160000001600000016", 
13965=>X"00000016000000160000001600000016", 13966=>X"00000016000000160000001600000016", 13967=>X"00000016000000160000001600000016", 13968=>X"00000016000000160000001600000016", 13969=>X"00000016000000160000001600000016", 
13970=>X"00000016000000160000001600000016", 13971=>X"00000016000000160000001600000016", 13972=>X"00000016000000160000001600000016", 13973=>X"00000016000000160000001600000016", 13974=>X"00000016000000160000001600000016", 
13975=>X"00000016000000160000001600000016", 13976=>X"00000016000000160000001600000016", 13977=>X"00000016000000160000001600000016", 13978=>X"00000016000000160000001600000016", 13979=>X"00000016000000160000001600000016", 
13980=>X"00000016000000160000001600000016", 13981=>X"00000016000000160000001600000016", 13982=>X"00000016000000160000001600000016", 13983=>X"00000016000000160000001600000016", 13984=>X"00000016000000160000001600000016", 
13985=>X"00000016000000160000001600000016", 13986=>X"00000016000000160000001600000016", 13987=>X"00000016000000160000001600000016", 13988=>X"00000016000000160000001600000016", 13989=>X"00000016000000160000001600000016", 
13990=>X"00000016000000160000001600000016", 13991=>X"00000016000000160000001600000016", 13992=>X"00000016000000160000001600000016", 13993=>X"00000016000000160000001600000016", 13994=>X"00000016000000160000001600000016", 
13995=>X"00000016000000160000001600000016", 13996=>X"00000016000000160000001600000016", 13997=>X"00000016000000160000001600000016", 13998=>X"00000016000000160000001600000016", 13999=>X"00000016000000160000001600000016", 
14000=>X"00000016000000160000001600000016", 14001=>X"00000016000000160000001600000016", 14002=>X"00000016000000160000001600000016", 14003=>X"00000016000000160000001600000016", 14004=>X"00000016000000160000001600000016", 
14005=>X"00000016000000160000001600000016", 14006=>X"00000016000000160000001600000016", 14007=>X"00000016000000160000001600000016", 14008=>X"00000016000000160000001600000016", 14009=>X"00000016000000160000001600000016", 
14010=>X"00000016000000160000001600000016", 14011=>X"00000016000000160000001600000016", 14012=>X"00000016000000160000001600000016", 14013=>X"00000016000000160000001600000016", 14014=>X"00000016000000160000001600000016", 
14015=>X"00000016000000160000001600000016", 14016=>X"00000016000000160000001600000016", 14017=>X"00000016000000160000001600000016", 14018=>X"00000016000000160000001600000016", 14019=>X"00000016000000160000001600000016", 
14020=>X"00000016000000160000001600000016", 14021=>X"00000016000000160000001600000016", 14022=>X"00000016000000160000001600000016", 14023=>X"00000016000000160000001600000016", 14024=>X"00000016000000160000001600000016", 
14025=>X"00000016000000160000001600000016", 14026=>X"00000016000000160000001600000016", 14027=>X"00000016000000160000001600000016", 14028=>X"00000016000000160000001600000016", 14029=>X"00000016000000160000001600000016", 
14030=>X"00000016000000160000001600000016", 14031=>X"00000016000000160000001600000016", 14032=>X"00000016000000160000001600000016", 14033=>X"00000016000000160000001600000016", 14034=>X"00000016000000160000001600000016", 
14035=>X"00000016000000160000001600000016", 14036=>X"00000016000000160000001600000016", 14037=>X"00000016000000160000001600000016", 14038=>X"00000016000000160000001600000016", 14039=>X"00000016000000160000001600000016", 
14040=>X"00000016000000160000001600000016", 14041=>X"00000016000000160000001600000016", 14042=>X"00000016000000160000001600000016", 14043=>X"00000016000000160000001600000016", 14044=>X"00000016000000160000001600000016", 
14045=>X"00000016000000160000001600000016", 14046=>X"00000016000000160000001600000016", 14047=>X"00000016000000160000001600000016", 14048=>X"00000016000000160000001600000016", 14049=>X"00000016000000160000001600000016", 
14050=>X"00000016000000160000001600000016", 14051=>X"00000016000000160000001600000016", 14052=>X"00000016000000160000001600000016", 14053=>X"00000016000000160000001600000016", 14054=>X"00000016000000160000001600000016", 
14055=>X"00000016000000160000001600000016", 14056=>X"00000016000000160000001600000016", 14057=>X"00000016000000160000001600000016", 14058=>X"00000016000000160000001600000016", 14059=>X"00000016000000160000001600000016", 
14060=>X"00000016000000160000001600000016", 14061=>X"00000016000000160000001600000016", 14062=>X"00000015000000150000001600000016", 14063=>X"00000015000000150000001500000015", 14064=>X"00000015000000150000001500000015", 
14065=>X"00000015000000150000001500000015", 14066=>X"00000015000000150000001500000015", 14067=>X"00000015000000150000001500000015", 14068=>X"00000015000000150000001500000015", 14069=>X"00000015000000150000001500000015", 
14070=>X"00000015000000150000001500000015", 14071=>X"00000015000000150000001500000015", 14072=>X"00000015000000150000001500000015", 14073=>X"00000015000000150000001500000015", 14074=>X"00000015000000150000001500000015", 
14075=>X"00000015000000150000001500000015", 14076=>X"00000015000000150000001500000015", 14077=>X"00000015000000150000001500000015", 14078=>X"00000015000000150000001500000015", 14079=>X"00000015000000150000001500000015", 
14080=>X"00000015000000150000001500000015", 14081=>X"00000015000000150000001500000015", 14082=>X"00000015000000150000001500000015", 14083=>X"00000015000000150000001500000015", 14084=>X"00000015000000150000001500000015", 
14085=>X"00000015000000150000001500000015", 14086=>X"00000015000000150000001500000015", 14087=>X"00000015000000150000001500000015", 14088=>X"00000015000000150000001500000015", 14089=>X"00000015000000150000001500000015", 
14090=>X"00000015000000150000001500000015", 14091=>X"00000015000000150000001500000015", 14092=>X"00000015000000150000001500000015", 14093=>X"00000015000000150000001500000015", 14094=>X"00000015000000150000001500000015", 
14095=>X"00000015000000150000001500000015", 14096=>X"00000015000000150000001500000015", 14097=>X"00000015000000150000001500000015", 14098=>X"00000015000000150000001500000015", 14099=>X"00000015000000150000001500000015", 
14100=>X"00000015000000150000001500000015", 14101=>X"00000015000000150000001500000015", 14102=>X"00000015000000150000001500000015", 14103=>X"00000015000000150000001500000015", 14104=>X"00000015000000150000001500000015", 
14105=>X"00000015000000150000001500000015", 14106=>X"00000015000000150000001500000015", 14107=>X"00000015000000150000001500000015", 14108=>X"00000015000000150000001500000015", 14109=>X"00000015000000150000001500000015", 
14110=>X"00000015000000150000001500000015", 14111=>X"00000015000000150000001500000015", 14112=>X"00000015000000150000001500000015", 14113=>X"00000015000000150000001500000015", 14114=>X"00000015000000150000001500000015", 
14115=>X"00000015000000150000001500000015", 14116=>X"00000015000000150000001500000015", 14117=>X"00000015000000150000001500000015", 14118=>X"00000015000000150000001500000015", 14119=>X"00000015000000150000001500000015", 
14120=>X"00000015000000150000001500000015", 14121=>X"00000015000000150000001500000015", 14122=>X"00000015000000150000001500000015", 14123=>X"00000015000000150000001500000015", 14124=>X"00000015000000150000001500000015", 
14125=>X"00000015000000150000001500000015", 14126=>X"00000015000000150000001500000015", 14127=>X"00000015000000150000001500000015", 14128=>X"00000015000000150000001500000015", 14129=>X"00000015000000150000001500000015", 
14130=>X"00000015000000150000001500000015", 14131=>X"00000015000000150000001500000015", 14132=>X"00000015000000150000001500000015", 14133=>X"00000015000000150000001500000015", 14134=>X"00000015000000150000001500000015", 
14135=>X"00000015000000150000001500000015", 14136=>X"00000015000000150000001500000015", 14137=>X"00000015000000150000001500000015", 14138=>X"00000015000000150000001500000015", 14139=>X"00000015000000150000001500000015", 
14140=>X"00000015000000150000001500000015", 14141=>X"00000015000000150000001500000015", 14142=>X"00000015000000150000001500000015", 14143=>X"00000015000000150000001500000015", 14144=>X"00000015000000150000001500000015", 
14145=>X"00000015000000150000001500000015", 14146=>X"00000015000000150000001500000015", 14147=>X"00000015000000150000001500000015", 14148=>X"00000015000000150000001500000015", 14149=>X"00000015000000150000001500000015", 
14150=>X"00000015000000150000001500000015", 14151=>X"00000015000000150000001500000015", 14152=>X"00000015000000150000001500000015", 14153=>X"00000015000000150000001500000015", 14154=>X"00000015000000150000001500000015", 
14155=>X"00000015000000150000001500000015", 14156=>X"00000015000000150000001500000015", 14157=>X"00000015000000150000001500000015", 14158=>X"00000015000000150000001500000015", 14159=>X"00000015000000150000001500000015", 
14160=>X"00000015000000150000001500000015", 14161=>X"00000015000000150000001500000015", 14162=>X"00000015000000150000001500000015", 14163=>X"00000015000000150000001500000015", 14164=>X"00000015000000150000001500000015", 
14165=>X"00000015000000150000001500000015", 14166=>X"00000015000000150000001500000015", 14167=>X"00000015000000150000001500000015", 14168=>X"00000015000000150000001500000015", 14169=>X"00000015000000150000001500000015", 
14170=>X"00000015000000150000001500000015", 14171=>X"00000015000000150000001500000015", 14172=>X"00000015000000150000001500000015", 14173=>X"00000015000000150000001500000015", 14174=>X"00000015000000150000001500000015", 
14175=>X"00000015000000150000001500000015", 14176=>X"00000015000000150000001500000015", 14177=>X"00000015000000150000001500000015", 14178=>X"00000015000000150000001500000015", 14179=>X"00000015000000150000001500000015", 
14180=>X"00000015000000150000001500000015", 14181=>X"00000015000000150000001500000015", 14182=>X"00000015000000150000001500000015", 14183=>X"00000015000000150000001500000015", 14184=>X"00000015000000150000001500000015", 
14185=>X"00000015000000150000001500000015", 14186=>X"00000015000000150000001500000015", 14187=>X"00000015000000150000001500000015", 14188=>X"00000015000000150000001500000015", 14189=>X"00000015000000150000001500000015", 
14190=>X"00000015000000150000001500000015", 14191=>X"00000015000000150000001500000015", 14192=>X"00000015000000150000001500000015", 14193=>X"00000015000000150000001500000015", 14194=>X"00000015000000150000001500000015", 
14195=>X"00000015000000150000001500000015", 14196=>X"00000015000000150000001500000015", 14197=>X"00000015000000150000001500000015", 14198=>X"00000015000000150000001500000015", 14199=>X"00000015000000150000001500000015", 
14200=>X"00000015000000150000001500000015", 14201=>X"00000015000000150000001500000015", 14202=>X"00000015000000150000001500000015", 14203=>X"00000015000000150000001500000015", 14204=>X"00000015000000150000001500000015", 
14205=>X"00000015000000150000001500000015", 14206=>X"00000015000000150000001500000015", 14207=>X"00000015000000150000001500000015", 14208=>X"00000015000000150000001500000015", 14209=>X"00000015000000150000001500000015", 
14210=>X"00000015000000150000001500000015", 14211=>X"00000015000000150000001500000015", 14212=>X"00000015000000150000001500000015", 14213=>X"00000015000000150000001500000015", 14214=>X"00000015000000150000001500000015", 
14215=>X"00000015000000150000001500000015", 14216=>X"00000015000000150000001500000015", 14217=>X"00000015000000150000001500000015", 14218=>X"00000015000000150000001500000015", 14219=>X"00000015000000150000001500000015", 
14220=>X"00000015000000150000001500000015", 14221=>X"00000015000000150000001500000015", 14222=>X"00000015000000150000001500000015", 14223=>X"00000015000000150000001500000015", 14224=>X"00000015000000150000001500000015", 
14225=>X"00000015000000150000001500000015", 14226=>X"00000015000000150000001500000015", 14227=>X"00000015000000150000001500000015", 14228=>X"00000015000000150000001500000015", 14229=>X"00000015000000150000001500000015", 
14230=>X"00000015000000150000001500000015", 14231=>X"00000015000000150000001500000015", 14232=>X"00000015000000150000001500000015", 14233=>X"00000015000000150000001500000015", 14234=>X"00000015000000150000001500000015", 
14235=>X"00000015000000150000001500000015", 14236=>X"00000015000000150000001500000015", 14237=>X"00000015000000150000001500000015", 14238=>X"00000015000000150000001500000015", 14239=>X"00000015000000150000001500000015", 
14240=>X"00000015000000150000001500000015", 14241=>X"00000015000000150000001500000015", 14242=>X"00000015000000150000001500000015", 14243=>X"00000015000000150000001500000015", 14244=>X"00000015000000150000001500000015", 
14245=>X"00000015000000150000001500000015", 14246=>X"00000015000000150000001500000015", 14247=>X"00000015000000150000001500000015", 14248=>X"00000015000000150000001500000015", 14249=>X"00000015000000150000001500000015", 
14250=>X"00000015000000150000001500000015", 14251=>X"00000015000000150000001500000015", 14252=>X"00000015000000150000001500000015", 14253=>X"00000015000000150000001500000015", 14254=>X"00000015000000150000001500000015", 
14255=>X"00000015000000150000001500000015", 14256=>X"00000015000000150000001500000015", 14257=>X"00000015000000150000001500000015", 14258=>X"00000015000000150000001500000015", 14259=>X"00000015000000150000001500000015", 
14260=>X"00000015000000150000001500000015", 14261=>X"00000015000000150000001500000015", 14262=>X"00000015000000150000001500000015", 14263=>X"00000015000000150000001500000015", 14264=>X"00000015000000150000001500000015", 
14265=>X"00000015000000150000001500000015", 14266=>X"00000015000000150000001500000015", 14267=>X"00000015000000150000001500000015", 14268=>X"00000015000000150000001500000015", 14269=>X"00000015000000150000001500000015", 
14270=>X"00000015000000150000001500000015", 14271=>X"00000015000000150000001500000015", 14272=>X"00000015000000150000001500000015", 14273=>X"00000015000000150000001500000015", 14274=>X"00000015000000150000001500000015", 
14275=>X"00000015000000150000001500000015", 14276=>X"00000015000000150000001500000015", 14277=>X"00000015000000150000001500000015", 14278=>X"00000015000000150000001500000015", 14279=>X"00000015000000150000001500000015", 
14280=>X"00000015000000150000001500000015", 14281=>X"00000015000000150000001500000015", 14282=>X"00000015000000150000001500000015", 14283=>X"00000015000000150000001500000015", 14284=>X"00000015000000150000001500000015", 
14285=>X"00000015000000150000001500000015", 14286=>X"00000015000000150000001500000015", 14287=>X"00000015000000150000001500000015", 14288=>X"00000015000000150000001500000015", 14289=>X"00000015000000150000001500000015", 
14290=>X"00000015000000150000001500000015", 14291=>X"00000015000000150000001500000015", 14292=>X"00000015000000150000001500000015", 14293=>X"00000015000000150000001500000015", 14294=>X"00000015000000150000001500000015", 
14295=>X"00000015000000150000001500000015", 14296=>X"00000015000000150000001500000015", 14297=>X"00000015000000150000001500000015", 14298=>X"00000015000000150000001500000015", 14299=>X"00000015000000150000001500000015", 
14300=>X"00000015000000150000001500000015", 14301=>X"00000015000000150000001500000015", 14302=>X"00000015000000150000001500000015", 14303=>X"00000015000000150000001500000015", 14304=>X"00000015000000150000001500000015", 
14305=>X"00000015000000150000001500000015", 14306=>X"00000015000000150000001500000015", 14307=>X"00000015000000150000001500000015", 14308=>X"00000015000000150000001500000015", 14309=>X"00000015000000150000001500000015", 
14310=>X"00000015000000150000001500000015", 14311=>X"00000015000000150000001500000015", 14312=>X"00000015000000150000001500000015", 14313=>X"00000015000000150000001500000015", 14314=>X"00000015000000150000001500000015", 
14315=>X"00000015000000150000001500000015", 14316=>X"00000015000000150000001500000015", 14317=>X"00000015000000150000001500000015", 14318=>X"00000015000000150000001500000015", 14319=>X"00000015000000150000001500000015", 
14320=>X"00000015000000150000001500000015", 14321=>X"00000015000000150000001500000015", 14322=>X"00000015000000150000001500000015", 14323=>X"00000015000000150000001500000015", 14324=>X"00000015000000150000001500000015", 
14325=>X"00000015000000150000001500000015", 14326=>X"00000015000000150000001500000015", 14327=>X"00000015000000150000001500000015", 14328=>X"00000015000000150000001500000015", 14329=>X"00000015000000150000001500000015", 
14330=>X"00000015000000150000001500000015", 14331=>X"00000015000000150000001500000015", 14332=>X"00000015000000150000001500000015", 14333=>X"00000015000000150000001500000015", 14334=>X"00000015000000150000001500000015", 
14335=>X"00000015000000150000001500000015", 14336=>X"00000015000000150000001500000015", 14337=>X"00000015000000150000001500000015", 14338=>X"00000015000000150000001500000015", 14339=>X"00000015000000150000001500000015", 
14340=>X"00000015000000150000001500000015", 14341=>X"00000015000000150000001500000015", 14342=>X"00000015000000150000001500000015", 14343=>X"00000015000000150000001500000015", 14344=>X"00000015000000150000001500000015", 
14345=>X"00000015000000150000001500000015", 14346=>X"00000015000000150000001500000015", 14347=>X"00000015000000150000001500000015", 14348=>X"00000015000000150000001500000015", 14349=>X"00000015000000150000001500000015", 
14350=>X"00000015000000150000001500000015", 14351=>X"00000015000000150000001500000015", 14352=>X"00000015000000150000001500000015", 14353=>X"00000015000000150000001500000015", 14354=>X"00000015000000150000001500000015", 
14355=>X"00000015000000150000001500000015", 14356=>X"00000015000000150000001500000015", 14357=>X"00000015000000150000001500000015", 14358=>X"00000015000000150000001500000015", 14359=>X"00000015000000150000001500000015", 
14360=>X"00000015000000150000001500000015", 14361=>X"00000015000000150000001500000015", 14362=>X"00000015000000150000001500000015", 14363=>X"00000015000000150000001500000015", 14364=>X"00000015000000150000001500000015", 
14365=>X"00000015000000150000001500000015", 14366=>X"00000015000000150000001500000015", 14367=>X"00000015000000150000001500000015", 14368=>X"00000015000000150000001500000015", 14369=>X"00000015000000150000001500000015", 
14370=>X"00000015000000150000001500000015", 14371=>X"00000015000000150000001500000015", 14372=>X"00000015000000150000001500000015", 14373=>X"00000015000000150000001500000015", 14374=>X"00000015000000150000001500000015", 
14375=>X"00000015000000150000001500000015", 14376=>X"00000015000000150000001500000015", 14377=>X"00000015000000150000001500000015", 14378=>X"00000015000000150000001500000015", 14379=>X"00000015000000150000001500000015", 
14380=>X"00000015000000150000001500000015", 14381=>X"00000015000000150000001500000015", 14382=>X"00000015000000150000001500000015", 14383=>X"00000015000000150000001500000015", 14384=>X"00000015000000150000001500000015", 
14385=>X"00000015000000150000001500000015", 14386=>X"00000015000000150000001500000015", 14387=>X"00000015000000150000001500000015", 14388=>X"00000015000000150000001500000015", 14389=>X"00000015000000150000001500000015", 
14390=>X"00000015000000150000001500000015", 14391=>X"00000015000000150000001500000015", 14392=>X"00000015000000150000001500000015", 14393=>X"00000015000000150000001500000015", 14394=>X"00000015000000150000001500000015", 
14395=>X"00000015000000150000001500000015", 14396=>X"00000015000000150000001500000015", 14397=>X"00000015000000150000001500000015", 14398=>X"00000015000000150000001500000015", 14399=>X"00000015000000150000001500000015", 
14400=>X"00000015000000150000001500000015", 14401=>X"00000015000000150000001500000015", 14402=>X"00000015000000150000001500000015", 14403=>X"00000015000000150000001500000015", 14404=>X"00000015000000150000001500000015", 
14405=>X"00000015000000150000001500000015", 14406=>X"00000015000000150000001500000015", 14407=>X"00000015000000150000001500000015", 14408=>X"00000015000000150000001500000015", 14409=>X"00000015000000150000001500000015", 
14410=>X"00000015000000150000001500000015", 14411=>X"00000015000000150000001500000015", 14412=>X"00000015000000150000001500000015", 14413=>X"00000015000000150000001500000015", 14414=>X"00000015000000150000001500000015", 
14415=>X"00000015000000150000001500000015", 14416=>X"00000015000000150000001500000015", 14417=>X"00000015000000150000001500000015", 14418=>X"00000015000000150000001500000015", 14419=>X"00000015000000150000001500000015", 
14420=>X"00000015000000150000001500000015", 14421=>X"00000015000000150000001500000015", 14422=>X"00000015000000150000001500000015", 14423=>X"00000015000000150000001500000015", 14424=>X"00000015000000150000001500000015", 
14425=>X"00000015000000150000001500000015", 14426=>X"00000015000000150000001500000015", 14427=>X"00000015000000150000001500000015", 14428=>X"00000015000000150000001500000015", 14429=>X"00000015000000150000001500000015", 
14430=>X"00000015000000150000001500000015", 14431=>X"00000015000000150000001500000015", 14432=>X"00000015000000150000001500000015", 14433=>X"00000015000000150000001500000015", 14434=>X"00000015000000150000001500000015", 
14435=>X"00000015000000150000001500000015", 14436=>X"00000015000000150000001500000015", 14437=>X"00000015000000150000001500000015", 14438=>X"00000015000000150000001500000015", 14439=>X"00000015000000150000001500000015", 
14440=>X"00000015000000150000001500000015", 14441=>X"00000015000000150000001500000015", 14442=>X"00000015000000150000001500000015", 14443=>X"00000015000000150000001500000015", 14444=>X"00000015000000150000001500000015", 
14445=>X"00000015000000150000001500000015", 14446=>X"00000015000000150000001500000015", 14447=>X"00000015000000150000001500000015", 14448=>X"00000015000000150000001500000015", 14449=>X"00000015000000150000001500000015", 
14450=>X"00000015000000150000001500000015", 14451=>X"00000015000000150000001500000015", 14452=>X"00000015000000150000001500000015", 14453=>X"00000015000000150000001500000015", 14454=>X"00000015000000150000001500000015", 
14455=>X"00000015000000150000001500000015", 14456=>X"00000015000000150000001500000015", 14457=>X"00000015000000150000001500000015", 14458=>X"00000015000000150000001500000015", 14459=>X"00000015000000150000001500000015", 
14460=>X"00000015000000150000001500000015", 14461=>X"00000015000000150000001500000015", 14462=>X"00000015000000150000001500000015", 14463=>X"00000015000000150000001500000015", 14464=>X"00000015000000150000001500000015", 
14465=>X"00000015000000150000001500000015", 14466=>X"00000015000000150000001500000015", 14467=>X"00000015000000150000001500000015", 14468=>X"00000015000000150000001500000015", 14469=>X"00000015000000150000001500000015", 
14470=>X"00000015000000150000001500000015", 14471=>X"00000015000000150000001500000015", 14472=>X"00000015000000150000001500000015", 14473=>X"00000015000000150000001500000015", 14474=>X"00000015000000150000001500000015", 
14475=>X"00000015000000150000001500000015", 14476=>X"00000015000000150000001500000015", 14477=>X"00000015000000150000001500000015", 14478=>X"00000015000000150000001500000015", 14479=>X"00000015000000150000001500000015", 
14480=>X"00000015000000150000001500000015", 14481=>X"00000015000000150000001500000015", 14482=>X"00000015000000150000001500000015", 14483=>X"00000015000000150000001500000015", 14484=>X"00000015000000150000001500000015", 
14485=>X"00000015000000150000001500000015", 14486=>X"00000015000000150000001500000015", 14487=>X"00000015000000150000001500000015", 14488=>X"00000015000000150000001500000015", 14489=>X"00000015000000150000001500000015", 
14490=>X"00000015000000150000001500000015", 14491=>X"00000015000000150000001500000015", 14492=>X"00000015000000150000001500000015", 14493=>X"00000015000000150000001500000015", 14494=>X"00000015000000150000001500000015", 
14495=>X"00000015000000150000001500000015", 14496=>X"00000015000000150000001500000015", 14497=>X"00000015000000150000001500000015", 14498=>X"00000015000000150000001500000015", 14499=>X"00000015000000150000001500000015", 
14500=>X"00000015000000150000001500000015", 14501=>X"00000015000000150000001500000015", 14502=>X"00000015000000150000001500000015", 14503=>X"00000015000000150000001500000015", 14504=>X"00000015000000150000001500000015", 
14505=>X"00000015000000150000001500000015", 14506=>X"00000015000000150000001500000015", 14507=>X"00000015000000150000001500000015", 14508=>X"00000015000000150000001500000015", 14509=>X"00000015000000150000001500000015", 
14510=>X"00000015000000150000001500000015", 14511=>X"00000015000000150000001500000015", 14512=>X"00000015000000150000001500000015", 14513=>X"00000015000000150000001500000015", 14514=>X"00000015000000150000001500000015", 
14515=>X"00000015000000150000001500000015", 14516=>X"00000015000000150000001500000015", 14517=>X"00000015000000150000001500000015", 14518=>X"00000015000000150000001500000015", 14519=>X"00000015000000150000001500000015", 
14520=>X"00000015000000150000001500000015", 14521=>X"00000015000000150000001500000015", 14522=>X"00000015000000150000001500000015", 14523=>X"00000015000000150000001500000015", 14524=>X"00000015000000150000001500000015", 
14525=>X"00000015000000150000001500000015", 14526=>X"00000015000000150000001500000015", 14527=>X"00000015000000150000001500000015", 14528=>X"00000015000000150000001500000015", 14529=>X"00000015000000150000001500000015", 
14530=>X"00000015000000150000001500000015", 14531=>X"00000015000000150000001500000015", 14532=>X"00000015000000150000001500000015", 14533=>X"00000015000000150000001500000015", 14534=>X"00000015000000150000001500000015", 
14535=>X"00000015000000150000001500000015", 14536=>X"00000015000000150000001500000015", 14537=>X"00000015000000150000001500000015", 14538=>X"00000015000000150000001500000015", 14539=>X"00000015000000150000001500000015", 
14540=>X"00000015000000150000001500000015", 14541=>X"00000015000000150000001500000015", 14542=>X"00000015000000150000001500000015", 14543=>X"00000015000000150000001500000015", 14544=>X"00000015000000150000001500000015", 
14545=>X"00000015000000150000001500000015", 14546=>X"00000015000000150000001500000015", 14547=>X"00000015000000150000001500000015", 14548=>X"00000015000000150000001500000015", 14549=>X"00000015000000150000001500000015", 
14550=>X"00000015000000150000001500000015", 14551=>X"00000015000000150000001500000015", 14552=>X"00000015000000150000001500000015", 14553=>X"00000015000000150000001500000015", 14554=>X"00000015000000150000001500000015", 
14555=>X"00000015000000150000001500000015", 14556=>X"00000015000000150000001500000015", 14557=>X"00000015000000150000001500000015", 14558=>X"00000015000000150000001500000015", 14559=>X"00000015000000150000001500000015", 
14560=>X"00000015000000150000001500000015", 14561=>X"00000015000000150000001500000015", 14562=>X"00000015000000150000001500000015", 14563=>X"00000015000000150000001500000015", 14564=>X"00000015000000150000001500000015", 
14565=>X"00000015000000150000001500000015", 14566=>X"00000015000000150000001500000015", 14567=>X"00000015000000150000001500000015", 14568=>X"00000015000000150000001500000015", 14569=>X"00000015000000150000001500000015", 
14570=>X"00000015000000150000001500000015", 14571=>X"00000015000000150000001500000015", 14572=>X"00000015000000150000001500000015", 14573=>X"00000015000000150000001500000015", 14574=>X"00000015000000150000001500000015", 
14575=>X"00000015000000150000001500000015", 14576=>X"00000015000000150000001500000015", 14577=>X"00000015000000150000001500000015", 14578=>X"00000015000000150000001500000015", 14579=>X"00000015000000150000001500000015", 
14580=>X"00000015000000150000001500000015", 14581=>X"00000015000000150000001500000015", 14582=>X"00000015000000150000001500000015", 14583=>X"00000015000000150000001500000015", 14584=>X"00000015000000150000001500000015", 
14585=>X"00000015000000150000001500000015", 14586=>X"00000015000000150000001500000015", 14587=>X"00000015000000150000001500000015", 14588=>X"00000015000000150000001500000015", 14589=>X"00000015000000150000001500000015", 
14590=>X"00000015000000150000001500000015", 14591=>X"00000015000000150000001500000015", 14592=>X"00000015000000150000001500000015", 14593=>X"00000015000000150000001500000015", 14594=>X"00000015000000150000001500000015", 
14595=>X"00000015000000150000001500000015", 14596=>X"00000015000000150000001500000015", 14597=>X"00000015000000150000001500000015", 14598=>X"00000015000000150000001500000015", 14599=>X"00000015000000150000001500000015", 
14600=>X"00000015000000150000001500000015", 14601=>X"00000015000000150000001500000015", 14602=>X"00000015000000150000001500000015", 14603=>X"00000015000000150000001500000015", 14604=>X"00000015000000150000001500000015", 
14605=>X"00000015000000150000001500000015", 14606=>X"00000015000000150000001500000015", 14607=>X"00000015000000150000001500000015", 14608=>X"00000015000000150000001500000015", 14609=>X"00000015000000150000001500000015", 
14610=>X"00000015000000150000001500000015", 14611=>X"00000015000000150000001500000015", 14612=>X"00000015000000150000001500000015", 14613=>X"00000015000000150000001500000015", 14614=>X"00000015000000150000001500000015", 
14615=>X"00000015000000150000001500000015", 14616=>X"00000015000000150000001500000015", 14617=>X"00000015000000150000001500000015", 14618=>X"00000015000000150000001500000015", 14619=>X"00000015000000150000001500000015", 
14620=>X"00000015000000150000001500000015", 14621=>X"00000015000000150000001500000015", 14622=>X"00000015000000150000001500000015", 14623=>X"00000015000000150000001500000015", 14624=>X"00000015000000150000001500000015", 
14625=>X"00000015000000150000001500000015", 14626=>X"00000015000000150000001500000015", 14627=>X"00000015000000150000001500000015", 14628=>X"00000015000000150000001500000015", 14629=>X"00000015000000150000001500000015", 
14630=>X"00000015000000150000001500000015", 14631=>X"00000015000000150000001500000015", 14632=>X"00000015000000150000001500000015", 14633=>X"00000015000000150000001500000015", 14634=>X"00000015000000150000001500000015", 
14635=>X"00000015000000150000001500000015", 14636=>X"00000015000000150000001500000015", 14637=>X"00000015000000150000001500000015", 14638=>X"00000015000000150000001500000015", 14639=>X"00000015000000150000001500000015", 
14640=>X"00000015000000150000001500000015", 14641=>X"00000015000000150000001500000015", 14642=>X"00000015000000150000001500000015", 14643=>X"00000015000000150000001500000015", 14644=>X"00000015000000150000001500000015", 
14645=>X"00000015000000150000001500000015", 14646=>X"00000015000000150000001500000015", 14647=>X"00000015000000150000001500000015", 14648=>X"00000015000000150000001500000015", 14649=>X"00000015000000150000001500000015", 
14650=>X"00000015000000150000001500000015", 14651=>X"00000015000000150000001500000015", 14652=>X"00000015000000150000001500000015", 14653=>X"00000015000000150000001500000015", 14654=>X"00000015000000150000001500000015", 
14655=>X"00000015000000150000001500000015", 14656=>X"00000015000000150000001500000015", 14657=>X"00000014000000140000001500000015", 14658=>X"00000014000000140000001400000014", 14659=>X"00000014000000140000001400000014", 
14660=>X"00000014000000140000001400000014", 14661=>X"00000014000000140000001400000014", 14662=>X"00000014000000140000001400000014", 14663=>X"00000014000000140000001400000014", 14664=>X"00000014000000140000001400000014", 
14665=>X"00000014000000140000001400000014", 14666=>X"00000014000000140000001400000014", 14667=>X"00000014000000140000001400000014", 14668=>X"00000014000000140000001400000014", 14669=>X"00000014000000140000001400000014", 
14670=>X"00000014000000140000001400000014", 14671=>X"00000014000000140000001400000014", 14672=>X"00000014000000140000001400000014", 14673=>X"00000014000000140000001400000014", 14674=>X"00000014000000140000001400000014", 
14675=>X"00000014000000140000001400000014", 14676=>X"00000014000000140000001400000014", 14677=>X"00000014000000140000001400000014", 14678=>X"00000014000000140000001400000014", 14679=>X"00000014000000140000001400000014", 
14680=>X"00000014000000140000001400000014", 14681=>X"00000014000000140000001400000014", 14682=>X"00000014000000140000001400000014", 14683=>X"00000014000000140000001400000014", 14684=>X"00000014000000140000001400000014", 
14685=>X"00000014000000140000001400000014", 14686=>X"00000014000000140000001400000014", 14687=>X"00000014000000140000001400000014", 14688=>X"00000014000000140000001400000014", 14689=>X"00000014000000140000001400000014", 
14690=>X"00000014000000140000001400000014", 14691=>X"00000014000000140000001400000014", 14692=>X"00000014000000140000001400000014", 14693=>X"00000014000000140000001400000014", 14694=>X"00000014000000140000001400000014", 
14695=>X"00000014000000140000001400000014", 14696=>X"00000014000000140000001400000014", 14697=>X"00000014000000140000001400000014", 14698=>X"00000014000000140000001400000014", 14699=>X"00000014000000140000001400000014", 
14700=>X"00000014000000140000001400000014", 14701=>X"00000014000000140000001400000014", 14702=>X"00000014000000140000001400000014", 14703=>X"00000014000000140000001400000014", 14704=>X"00000014000000140000001400000014", 
14705=>X"00000014000000140000001400000014", 14706=>X"00000014000000140000001400000014", 14707=>X"00000014000000140000001400000014", 14708=>X"00000014000000140000001400000014", 14709=>X"00000014000000140000001400000014", 
14710=>X"00000014000000140000001400000014", 14711=>X"00000014000000140000001400000014", 14712=>X"00000014000000140000001400000014", 14713=>X"00000014000000140000001400000014", 14714=>X"00000014000000140000001400000014", 
14715=>X"00000014000000140000001400000014", 14716=>X"00000014000000140000001400000014", 14717=>X"00000014000000140000001400000014", 14718=>X"00000014000000140000001400000014", 14719=>X"00000014000000140000001400000014", 
14720=>X"00000014000000140000001400000014", 14721=>X"00000014000000140000001400000014", 14722=>X"00000014000000140000001400000014", 14723=>X"00000014000000140000001400000014", 14724=>X"00000014000000140000001400000014", 
14725=>X"00000014000000140000001400000014", 14726=>X"00000014000000140000001400000014", 14727=>X"00000014000000140000001400000014", 14728=>X"00000014000000140000001400000014", 14729=>X"00000014000000140000001400000014", 
14730=>X"00000014000000140000001400000014", 14731=>X"00000014000000140000001400000014", 14732=>X"00000014000000140000001400000014", 14733=>X"00000014000000140000001400000014", 14734=>X"00000014000000140000001400000014", 
14735=>X"00000014000000140000001400000014", 14736=>X"00000014000000140000001400000014", 14737=>X"00000014000000140000001400000014", 14738=>X"00000014000000140000001400000014", 14739=>X"00000014000000140000001400000014", 
14740=>X"00000014000000140000001400000014", 14741=>X"00000014000000140000001400000014", 14742=>X"00000014000000140000001400000014", 14743=>X"00000014000000140000001400000014", 14744=>X"00000014000000140000001400000014", 
14745=>X"00000014000000140000001400000014", 14746=>X"00000014000000140000001400000014", 14747=>X"00000014000000140000001400000014", 14748=>X"00000014000000140000001400000014", 14749=>X"00000014000000140000001400000014", 
14750=>X"00000014000000140000001400000014", 14751=>X"00000014000000140000001400000014", 14752=>X"00000014000000140000001400000014", 14753=>X"00000014000000140000001400000014", 14754=>X"00000014000000140000001400000014", 
14755=>X"00000014000000140000001400000014", 14756=>X"00000014000000140000001400000014", 14757=>X"00000014000000140000001400000014", 14758=>X"00000014000000140000001400000014", 14759=>X"00000014000000140000001400000014", 
14760=>X"00000014000000140000001400000014", 14761=>X"00000014000000140000001400000014", 14762=>X"00000014000000140000001400000014", 14763=>X"00000014000000140000001400000014", 14764=>X"00000014000000140000001400000014", 
14765=>X"00000014000000140000001400000014", 14766=>X"00000014000000140000001400000014", 14767=>X"00000014000000140000001400000014", 14768=>X"00000014000000140000001400000014", 14769=>X"00000014000000140000001400000014", 
14770=>X"00000014000000140000001400000014", 14771=>X"00000014000000140000001400000014", 14772=>X"00000014000000140000001400000014", 14773=>X"00000014000000140000001400000014", 14774=>X"00000014000000140000001400000014", 
14775=>X"00000014000000140000001400000014", 14776=>X"00000014000000140000001400000014", 14777=>X"00000014000000140000001400000014", 14778=>X"00000014000000140000001400000014", 14779=>X"00000014000000140000001400000014", 
14780=>X"00000014000000140000001400000014", 14781=>X"00000014000000140000001400000014", 14782=>X"00000014000000140000001400000014", 14783=>X"00000014000000140000001400000014", 14784=>X"00000014000000140000001400000014", 
14785=>X"00000014000000140000001400000014", 14786=>X"00000014000000140000001400000014", 14787=>X"00000014000000140000001400000014", 14788=>X"00000014000000140000001400000014", 14789=>X"00000014000000140000001400000014", 
14790=>X"00000014000000140000001400000014", 14791=>X"00000014000000140000001400000014", 14792=>X"00000014000000140000001400000014", 14793=>X"00000014000000140000001400000014", 14794=>X"00000014000000140000001400000014", 
14795=>X"00000014000000140000001400000014", 14796=>X"00000014000000140000001400000014", 14797=>X"00000014000000140000001400000014", 14798=>X"00000014000000140000001400000014", 14799=>X"00000014000000140000001400000014", 
14800=>X"00000014000000140000001400000014", 14801=>X"00000014000000140000001400000014", 14802=>X"00000014000000140000001400000014", 14803=>X"00000014000000140000001400000014", 14804=>X"00000014000000140000001400000014", 
14805=>X"00000014000000140000001400000014", 14806=>X"00000014000000140000001400000014", 14807=>X"00000014000000140000001400000014", 14808=>X"00000014000000140000001400000014", 14809=>X"00000014000000140000001400000014", 
14810=>X"00000014000000140000001400000014", 14811=>X"00000014000000140000001400000014", 14812=>X"00000014000000140000001400000014", 14813=>X"00000014000000140000001400000014", 14814=>X"00000014000000140000001400000014", 
14815=>X"00000014000000140000001400000014", 14816=>X"00000014000000140000001400000014", 14817=>X"00000014000000140000001400000014", 14818=>X"00000014000000140000001400000014", 14819=>X"00000014000000140000001400000014", 
14820=>X"00000014000000140000001400000014", 14821=>X"00000014000000140000001400000014", 14822=>X"00000014000000140000001400000014", 14823=>X"00000014000000140000001400000014", 14824=>X"00000014000000140000001400000014", 
14825=>X"00000014000000140000001400000014", 14826=>X"00000014000000140000001400000014", 14827=>X"00000014000000140000001400000014", 14828=>X"00000014000000140000001400000014", 14829=>X"00000014000000140000001400000014", 
14830=>X"00000014000000140000001400000014", 14831=>X"00000014000000140000001400000014", 14832=>X"00000014000000140000001400000014", 14833=>X"00000014000000140000001400000014", 14834=>X"00000014000000140000001400000014", 
14835=>X"00000014000000140000001400000014", 14836=>X"00000014000000140000001400000014", 14837=>X"00000014000000140000001400000014", 14838=>X"00000014000000140000001400000014", 14839=>X"00000014000000140000001400000014", 
14840=>X"00000014000000140000001400000014", 14841=>X"00000014000000140000001400000014", 14842=>X"00000014000000140000001400000014", 14843=>X"00000014000000140000001400000014", 14844=>X"00000014000000140000001400000014", 
14845=>X"00000014000000140000001400000014", 14846=>X"00000014000000140000001400000014", 14847=>X"00000014000000140000001400000014", 14848=>X"00000014000000140000001400000014", 14849=>X"00000014000000140000001400000014", 
14850=>X"00000014000000140000001400000014", 14851=>X"00000014000000140000001400000014", 14852=>X"00000014000000140000001400000014", 14853=>X"00000014000000140000001400000014", 14854=>X"00000014000000140000001400000014", 
14855=>X"00000014000000140000001400000014", 14856=>X"00000014000000140000001400000014", 14857=>X"00000014000000140000001400000014", 14858=>X"00000014000000140000001400000014", 14859=>X"00000014000000140000001400000014", 
14860=>X"00000014000000140000001400000014", 14861=>X"00000014000000140000001400000014", 14862=>X"00000014000000140000001400000014", 14863=>X"00000014000000140000001400000014", 14864=>X"00000014000000140000001400000014", 
14865=>X"00000014000000140000001400000014", 14866=>X"00000014000000140000001400000014", 14867=>X"00000014000000140000001400000014", 14868=>X"00000014000000140000001400000014", 14869=>X"00000014000000140000001400000014", 
14870=>X"00000014000000140000001400000014", 14871=>X"00000014000000140000001400000014", 14872=>X"00000014000000140000001400000014", 14873=>X"00000014000000140000001400000014", 14874=>X"00000014000000140000001400000014", 
14875=>X"00000014000000140000001400000014", 14876=>X"00000014000000140000001400000014", 14877=>X"00000014000000140000001400000014", 14878=>X"00000014000000140000001400000014", 14879=>X"00000014000000140000001400000014", 
14880=>X"00000014000000140000001400000014", 14881=>X"00000014000000140000001400000014", 14882=>X"00000014000000140000001400000014", 14883=>X"00000014000000140000001400000014", 14884=>X"00000014000000140000001400000014", 
14885=>X"00000014000000140000001400000014", 14886=>X"00000014000000140000001400000014", 14887=>X"00000014000000140000001400000014", 14888=>X"00000014000000140000001400000014", 14889=>X"00000014000000140000001400000014", 
14890=>X"00000014000000140000001400000014", 14891=>X"00000014000000140000001400000014", 14892=>X"00000014000000140000001400000014", 14893=>X"00000014000000140000001400000014", 14894=>X"00000014000000140000001400000014", 
14895=>X"00000014000000140000001400000014", 14896=>X"00000014000000140000001400000014", 14897=>X"00000014000000140000001400000014", 14898=>X"00000014000000140000001400000014", 14899=>X"00000014000000140000001400000014", 
14900=>X"00000014000000140000001400000014", 14901=>X"00000014000000140000001400000014", 14902=>X"00000014000000140000001400000014", 14903=>X"00000014000000140000001400000014", 14904=>X"00000014000000140000001400000014", 
14905=>X"00000014000000140000001400000014", 14906=>X"00000014000000140000001400000014", 14907=>X"00000014000000140000001400000014", 14908=>X"00000014000000140000001400000014", 14909=>X"00000014000000140000001400000014", 
14910=>X"00000014000000140000001400000014", 14911=>X"00000014000000140000001400000014", 14912=>X"00000014000000140000001400000014", 14913=>X"00000014000000140000001400000014", 14914=>X"00000014000000140000001400000014", 
14915=>X"00000014000000140000001400000014", 14916=>X"00000014000000140000001400000014", 14917=>X"00000014000000140000001400000014", 14918=>X"00000014000000140000001400000014", 14919=>X"00000014000000140000001400000014", 
14920=>X"00000014000000140000001400000014", 14921=>X"00000014000000140000001400000014", 14922=>X"00000014000000140000001400000014", 14923=>X"00000014000000140000001400000014", 14924=>X"00000014000000140000001400000014", 
14925=>X"00000014000000140000001400000014", 14926=>X"00000014000000140000001400000014", 14927=>X"00000014000000140000001400000014", 14928=>X"00000014000000140000001400000014", 14929=>X"00000014000000140000001400000014", 
14930=>X"00000014000000140000001400000014", 14931=>X"00000014000000140000001400000014", 14932=>X"00000014000000140000001400000014", 14933=>X"00000014000000140000001400000014", 14934=>X"00000014000000140000001400000014", 
14935=>X"00000014000000140000001400000014", 14936=>X"00000014000000140000001400000014", 14937=>X"00000014000000140000001400000014", 14938=>X"00000014000000140000001400000014", 14939=>X"00000014000000140000001400000014", 
14940=>X"00000014000000140000001400000014", 14941=>X"00000014000000140000001400000014", 14942=>X"00000014000000140000001400000014", 14943=>X"00000014000000140000001400000014", 14944=>X"00000014000000140000001400000014", 
14945=>X"00000014000000140000001400000014", 14946=>X"00000014000000140000001400000014", 14947=>X"00000014000000140000001400000014", 14948=>X"00000014000000140000001400000014", 14949=>X"00000014000000140000001400000014", 
14950=>X"00000014000000140000001400000014", 14951=>X"00000014000000140000001400000014", 14952=>X"00000014000000140000001400000014", 14953=>X"00000014000000140000001400000014", 14954=>X"00000014000000140000001400000014", 
14955=>X"00000014000000140000001400000014", 14956=>X"00000014000000140000001400000014", 14957=>X"00000014000000140000001400000014", 14958=>X"00000014000000140000001400000014", 14959=>X"00000014000000140000001400000014", 
14960=>X"00000014000000140000001400000014", 14961=>X"00000014000000140000001400000014", 14962=>X"00000014000000140000001400000014", 14963=>X"00000014000000140000001400000014", 14964=>X"00000014000000140000001400000014", 
14965=>X"00000014000000140000001400000014", 14966=>X"00000014000000140000001400000014", 14967=>X"00000014000000140000001400000014", 14968=>X"00000014000000140000001400000014", 14969=>X"00000014000000140000001400000014", 
14970=>X"00000014000000140000001400000014", 14971=>X"00000014000000140000001400000014", 14972=>X"00000014000000140000001400000014", 14973=>X"00000014000000140000001400000014", 14974=>X"00000014000000140000001400000014", 
14975=>X"00000014000000140000001400000014", 14976=>X"00000014000000140000001400000014", 14977=>X"00000014000000140000001400000014", 14978=>X"00000014000000140000001400000014", 14979=>X"00000014000000140000001400000014", 
14980=>X"00000014000000140000001400000014", 14981=>X"00000014000000140000001400000014", 14982=>X"00000014000000140000001400000014", 14983=>X"00000014000000140000001400000014", 14984=>X"00000014000000140000001400000014", 
14985=>X"00000014000000140000001400000014", 14986=>X"00000014000000140000001400000014", 14987=>X"00000014000000140000001400000014", 14988=>X"00000014000000140000001400000014", 14989=>X"00000014000000140000001400000014", 
14990=>X"00000014000000140000001400000014", 14991=>X"00000014000000140000001400000014", 14992=>X"00000014000000140000001400000014", 14993=>X"00000014000000140000001400000014", 14994=>X"00000014000000140000001400000014", 
14995=>X"00000014000000140000001400000014", 14996=>X"00000014000000140000001400000014", 14997=>X"00000014000000140000001400000014", 14998=>X"00000014000000140000001400000014", 14999=>X"00000014000000140000001400000014", 
15000=>X"00000014000000140000001400000014", 15001=>X"00000014000000140000001400000014", 15002=>X"00000014000000140000001400000014", 15003=>X"00000014000000140000001400000014", 15004=>X"00000014000000140000001400000014", 
15005=>X"00000014000000140000001400000014", 15006=>X"00000014000000140000001400000014", 15007=>X"00000014000000140000001400000014", 15008=>X"00000014000000140000001400000014", 15009=>X"00000014000000140000001400000014", 
15010=>X"00000014000000140000001400000014", 15011=>X"00000014000000140000001400000014", 15012=>X"00000014000000140000001400000014", 15013=>X"00000014000000140000001400000014", 15014=>X"00000014000000140000001400000014", 
15015=>X"00000014000000140000001400000014", 15016=>X"00000014000000140000001400000014", 15017=>X"00000014000000140000001400000014", 15018=>X"00000014000000140000001400000014", 15019=>X"00000014000000140000001400000014", 
15020=>X"00000014000000140000001400000014", 15021=>X"00000014000000140000001400000014", 15022=>X"00000014000000140000001400000014", 15023=>X"00000014000000140000001400000014", 15024=>X"00000014000000140000001400000014", 
15025=>X"00000014000000140000001400000014", 15026=>X"00000014000000140000001400000014", 15027=>X"00000014000000140000001400000014", 15028=>X"00000014000000140000001400000014", 15029=>X"00000014000000140000001400000014", 
15030=>X"00000014000000140000001400000014", 15031=>X"00000014000000140000001400000014", 15032=>X"00000014000000140000001400000014", 15033=>X"00000014000000140000001400000014", 15034=>X"00000014000000140000001400000014", 
15035=>X"00000014000000140000001400000014", 15036=>X"00000014000000140000001400000014", 15037=>X"00000014000000140000001400000014", 15038=>X"00000014000000140000001400000014", 15039=>X"00000014000000140000001400000014", 
15040=>X"00000014000000140000001400000014", 15041=>X"00000014000000140000001400000014", 15042=>X"00000014000000140000001400000014", 15043=>X"00000014000000140000001400000014", 15044=>X"00000014000000140000001400000014", 
15045=>X"00000014000000140000001400000014", 15046=>X"00000014000000140000001400000014", 15047=>X"00000014000000140000001400000014", 15048=>X"00000014000000140000001400000014", 15049=>X"00000014000000140000001400000014", 
15050=>X"00000014000000140000001400000014", 15051=>X"00000014000000140000001400000014", 15052=>X"00000014000000140000001400000014", 15053=>X"00000014000000140000001400000014", 15054=>X"00000014000000140000001400000014", 
15055=>X"00000014000000140000001400000014", 15056=>X"00000014000000140000001400000014", 15057=>X"00000014000000140000001400000014", 15058=>X"00000014000000140000001400000014", 15059=>X"00000014000000140000001400000014", 
15060=>X"00000014000000140000001400000014", 15061=>X"00000014000000140000001400000014", 15062=>X"00000014000000140000001400000014", 15063=>X"00000014000000140000001400000014", 15064=>X"00000014000000140000001400000014", 
15065=>X"00000014000000140000001400000014", 15066=>X"00000014000000140000001400000014", 15067=>X"00000014000000140000001400000014", 15068=>X"00000014000000140000001400000014", 15069=>X"00000014000000140000001400000014", 
15070=>X"00000014000000140000001400000014", 15071=>X"00000014000000140000001400000014", 15072=>X"00000014000000140000001400000014", 15073=>X"00000014000000140000001400000014", 15074=>X"00000014000000140000001400000014", 
15075=>X"00000014000000140000001400000014", 15076=>X"00000014000000140000001400000014", 15077=>X"00000014000000140000001400000014", 15078=>X"00000014000000140000001400000014", 15079=>X"00000014000000140000001400000014", 
15080=>X"00000014000000140000001400000014", 15081=>X"00000014000000140000001400000014", 15082=>X"00000014000000140000001400000014", 15083=>X"00000014000000140000001400000014", 15084=>X"00000014000000140000001400000014", 
15085=>X"00000014000000140000001400000014", 15086=>X"00000014000000140000001400000014", 15087=>X"00000014000000140000001400000014", 15088=>X"00000014000000140000001400000014", 15089=>X"00000014000000140000001400000014", 
15090=>X"00000014000000140000001400000014", 15091=>X"00000014000000140000001400000014", 15092=>X"00000014000000140000001400000014", 15093=>X"00000014000000140000001400000014", 15094=>X"00000014000000140000001400000014", 
15095=>X"00000014000000140000001400000014", 15096=>X"00000014000000140000001400000014", 15097=>X"00000014000000140000001400000014", 15098=>X"00000014000000140000001400000014", 15099=>X"00000014000000140000001400000014", 
15100=>X"00000014000000140000001400000014", 15101=>X"00000014000000140000001400000014", 15102=>X"00000014000000140000001400000014", 15103=>X"00000014000000140000001400000014", 15104=>X"00000014000000140000001400000014", 
15105=>X"00000014000000140000001400000014", 15106=>X"00000014000000140000001400000014", 15107=>X"00000014000000140000001400000014", 15108=>X"00000014000000140000001400000014", 15109=>X"00000014000000140000001400000014", 
15110=>X"00000014000000140000001400000014", 15111=>X"00000014000000140000001400000014", 15112=>X"00000014000000140000001400000014", 15113=>X"00000014000000140000001400000014", 15114=>X"00000014000000140000001400000014", 
15115=>X"00000014000000140000001400000014", 15116=>X"00000014000000140000001400000014", 15117=>X"00000014000000140000001400000014", 15118=>X"00000014000000140000001400000014", 15119=>X"00000014000000140000001400000014", 
15120=>X"00000014000000140000001400000014", 15121=>X"00000014000000140000001400000014", 15122=>X"00000014000000140000001400000014", 15123=>X"00000014000000140000001400000014", 15124=>X"00000014000000140000001400000014", 
15125=>X"00000014000000140000001400000014", 15126=>X"00000014000000140000001400000014", 15127=>X"00000014000000140000001400000014", 15128=>X"00000014000000140000001400000014", 15129=>X"00000014000000140000001400000014", 
15130=>X"00000014000000140000001400000014", 15131=>X"00000014000000140000001400000014", 15132=>X"00000014000000140000001400000014", 15133=>X"00000014000000140000001400000014", 15134=>X"00000014000000140000001400000014", 
15135=>X"00000014000000140000001400000014", 15136=>X"00000014000000140000001400000014", 15137=>X"00000014000000140000001400000014", 15138=>X"00000014000000140000001400000014", 15139=>X"00000014000000140000001400000014", 
15140=>X"00000014000000140000001400000014", 15141=>X"00000014000000140000001400000014", 15142=>X"00000014000000140000001400000014", 15143=>X"00000014000000140000001400000014", 15144=>X"00000014000000140000001400000014", 
15145=>X"00000014000000140000001400000014", 15146=>X"00000014000000140000001400000014", 15147=>X"00000014000000140000001400000014", 15148=>X"00000014000000140000001400000014", 15149=>X"00000014000000140000001400000014", 
15150=>X"00000014000000140000001400000014", 15151=>X"00000014000000140000001400000014", 15152=>X"00000014000000140000001400000014", 15153=>X"00000014000000140000001400000014", 15154=>X"00000014000000140000001400000014", 
15155=>X"00000014000000140000001400000014", 15156=>X"00000014000000140000001400000014", 15157=>X"00000014000000140000001400000014", 15158=>X"00000014000000140000001400000014", 15159=>X"00000014000000140000001400000014", 
15160=>X"00000014000000140000001400000014", 15161=>X"00000014000000140000001400000014", 15162=>X"00000014000000140000001400000014", 15163=>X"00000014000000140000001400000014", 15164=>X"00000014000000140000001400000014", 
15165=>X"00000014000000140000001400000014", 15166=>X"00000014000000140000001400000014", 15167=>X"00000014000000140000001400000014", 15168=>X"00000014000000140000001400000014", 15169=>X"00000014000000140000001400000014", 
15170=>X"00000014000000140000001400000014", 15171=>X"00000014000000140000001400000014", 15172=>X"00000014000000140000001400000014", 15173=>X"00000014000000140000001400000014", 15174=>X"00000014000000140000001400000014", 
15175=>X"00000014000000140000001400000014", 15176=>X"00000014000000140000001400000014", 15177=>X"00000014000000140000001400000014", 15178=>X"00000014000000140000001400000014", 15179=>X"00000014000000140000001400000014", 
15180=>X"00000014000000140000001400000014", 15181=>X"00000014000000140000001400000014", 15182=>X"00000014000000140000001400000014", 15183=>X"00000014000000140000001400000014", 15184=>X"00000014000000140000001400000014", 
15185=>X"00000014000000140000001400000014", 15186=>X"00000014000000140000001400000014", 15187=>X"00000014000000140000001400000014", 15188=>X"00000014000000140000001400000014", 15189=>X"00000014000000140000001400000014", 
15190=>X"00000014000000140000001400000014", 15191=>X"00000014000000140000001400000014", 15192=>X"00000014000000140000001400000014", 15193=>X"00000014000000140000001400000014", 15194=>X"00000014000000140000001400000014", 
15195=>X"00000014000000140000001400000014", 15196=>X"00000014000000140000001400000014", 15197=>X"00000014000000140000001400000014", 15198=>X"00000014000000140000001400000014", 15199=>X"00000014000000140000001400000014", 
15200=>X"00000014000000140000001400000014", 15201=>X"00000014000000140000001400000014", 15202=>X"00000014000000140000001400000014", 15203=>X"00000014000000140000001400000014", 15204=>X"00000014000000140000001400000014", 
15205=>X"00000014000000140000001400000014", 15206=>X"00000014000000140000001400000014", 15207=>X"00000014000000140000001400000014", 15208=>X"00000014000000140000001400000014", 15209=>X"00000014000000140000001400000014", 
15210=>X"00000014000000140000001400000014", 15211=>X"00000014000000140000001400000014", 15212=>X"00000014000000140000001400000014", 15213=>X"00000014000000140000001400000014", 15214=>X"00000014000000140000001400000014", 
15215=>X"00000014000000140000001400000014", 15216=>X"00000014000000140000001400000014", 15217=>X"00000014000000140000001400000014", 15218=>X"00000014000000140000001400000014", 15219=>X"00000014000000140000001400000014", 
15220=>X"00000014000000140000001400000014", 15221=>X"00000014000000140000001400000014", 15222=>X"00000014000000140000001400000014", 15223=>X"00000014000000140000001400000014", 15224=>X"00000014000000140000001400000014", 
15225=>X"00000014000000140000001400000014", 15226=>X"00000014000000140000001400000014", 15227=>X"00000014000000140000001400000014", 15228=>X"00000014000000140000001400000014", 15229=>X"00000014000000140000001400000014", 
15230=>X"00000014000000140000001400000014", 15231=>X"00000014000000140000001400000014", 15232=>X"00000014000000140000001400000014", 15233=>X"00000014000000140000001400000014", 15234=>X"00000014000000140000001400000014", 
15235=>X"00000014000000140000001400000014", 15236=>X"00000014000000140000001400000014", 15237=>X"00000014000000140000001400000014", 15238=>X"00000014000000140000001400000014", 15239=>X"00000014000000140000001400000014", 
15240=>X"00000014000000140000001400000014", 15241=>X"00000014000000140000001400000014", 15242=>X"00000014000000140000001400000014", 15243=>X"00000014000000140000001400000014", 15244=>X"00000014000000140000001400000014", 
15245=>X"00000014000000140000001400000014", 15246=>X"00000014000000140000001400000014", 15247=>X"00000014000000140000001400000014", 15248=>X"00000014000000140000001400000014", 15249=>X"00000014000000140000001400000014", 
15250=>X"00000014000000140000001400000014", 15251=>X"00000014000000140000001400000014", 15252=>X"00000014000000140000001400000014", 15253=>X"00000014000000140000001400000014", 15254=>X"00000014000000140000001400000014", 
15255=>X"00000014000000140000001400000014", 15256=>X"00000014000000140000001400000014", 15257=>X"00000014000000140000001400000014", 15258=>X"00000014000000140000001400000014", 15259=>X"00000014000000140000001400000014", 
15260=>X"00000014000000140000001400000014", 15261=>X"00000014000000140000001400000014", 15262=>X"00000014000000140000001400000014", 15263=>X"00000014000000140000001400000014", 15264=>X"00000014000000140000001400000014", 
15265=>X"00000014000000140000001400000014", 15266=>X"00000014000000140000001400000014", 15267=>X"00000014000000140000001400000014", 15268=>X"00000014000000140000001400000014", 15269=>X"00000014000000140000001400000014", 
15270=>X"00000014000000140000001400000014", 15271=>X"00000014000000140000001400000014", 15272=>X"00000014000000140000001400000014", 15273=>X"00000014000000140000001400000014", 15274=>X"00000014000000140000001400000014", 
15275=>X"00000014000000140000001400000014", 15276=>X"00000014000000140000001400000014", 15277=>X"00000014000000140000001400000014", 15278=>X"00000014000000140000001400000014", 15279=>X"00000014000000140000001400000014", 
15280=>X"00000014000000140000001400000014", 15281=>X"00000014000000140000001400000014", 15282=>X"00000014000000140000001400000014", 15283=>X"00000014000000140000001400000014", 15284=>X"00000014000000140000001400000014", 
15285=>X"00000014000000140000001400000014", 15286=>X"00000014000000140000001400000014", 15287=>X"00000014000000140000001400000014", 15288=>X"00000014000000140000001400000014", 15289=>X"00000014000000140000001400000014", 
15290=>X"00000014000000140000001400000014", 15291=>X"00000014000000140000001400000014", 15292=>X"00000014000000140000001400000014", 15293=>X"00000014000000140000001400000014", 15294=>X"00000014000000140000001400000014", 
15295=>X"00000014000000140000001400000014", 15296=>X"00000014000000140000001400000014", 15297=>X"00000014000000140000001400000014", 15298=>X"00000014000000140000001400000014", 15299=>X"00000014000000140000001400000014", 
15300=>X"00000014000000140000001400000014", 15301=>X"00000014000000140000001400000014", 15302=>X"00000014000000140000001400000014", 15303=>X"00000014000000140000001400000014", 15304=>X"00000014000000140000001400000014", 
15305=>X"00000014000000140000001400000014", 15306=>X"00000014000000140000001400000014", 15307=>X"00000014000000140000001400000014", 15308=>X"00000014000000140000001400000014", 15309=>X"00000014000000140000001400000014", 
15310=>X"00000014000000140000001400000014", 15311=>X"00000014000000140000001400000014", 15312=>X"00000014000000140000001400000014", 15313=>X"00000013000000130000001300000014", 15314=>X"00000013000000130000001300000013", 
15315=>X"00000013000000130000001300000013", 15316=>X"00000013000000130000001300000013", 15317=>X"00000013000000130000001300000013", 15318=>X"00000013000000130000001300000013", 15319=>X"00000013000000130000001300000013", 
15320=>X"00000013000000130000001300000013", 15321=>X"00000013000000130000001300000013", 15322=>X"00000013000000130000001300000013", 15323=>X"00000013000000130000001300000013", 15324=>X"00000013000000130000001300000013", 
15325=>X"00000013000000130000001300000013", 15326=>X"00000013000000130000001300000013", 15327=>X"00000013000000130000001300000013", 15328=>X"00000013000000130000001300000013", 15329=>X"00000013000000130000001300000013", 
15330=>X"00000013000000130000001300000013", 15331=>X"00000013000000130000001300000013", 15332=>X"00000013000000130000001300000013", 15333=>X"00000013000000130000001300000013", 15334=>X"00000013000000130000001300000013", 
15335=>X"00000013000000130000001300000013", 15336=>X"00000013000000130000001300000013", 15337=>X"00000013000000130000001300000013", 15338=>X"00000013000000130000001300000013", 15339=>X"00000013000000130000001300000013", 
15340=>X"00000013000000130000001300000013", 15341=>X"00000013000000130000001300000013", 15342=>X"00000013000000130000001300000013", 15343=>X"00000013000000130000001300000013", 15344=>X"00000013000000130000001300000013", 
15345=>X"00000013000000130000001300000013", 15346=>X"00000013000000130000001300000013", 15347=>X"00000013000000130000001300000013", 15348=>X"00000013000000130000001300000013", 15349=>X"00000013000000130000001300000013", 
15350=>X"00000013000000130000001300000013", 15351=>X"00000013000000130000001300000013", 15352=>X"00000013000000130000001300000013", 15353=>X"00000013000000130000001300000013", 15354=>X"00000013000000130000001300000013", 
15355=>X"00000013000000130000001300000013", 15356=>X"00000013000000130000001300000013", 15357=>X"00000013000000130000001300000013", 15358=>X"00000013000000130000001300000013", 15359=>X"00000013000000130000001300000013", 
15360=>X"00000013000000130000001300000013", 15361=>X"00000013000000130000001300000013", 15362=>X"00000013000000130000001300000013", 15363=>X"00000013000000130000001300000013", 15364=>X"00000013000000130000001300000013", 
15365=>X"00000013000000130000001300000013", 15366=>X"00000013000000130000001300000013", 15367=>X"00000013000000130000001300000013", 15368=>X"00000013000000130000001300000013", 15369=>X"00000013000000130000001300000013", 
15370=>X"00000013000000130000001300000013", 15371=>X"00000013000000130000001300000013", 15372=>X"00000013000000130000001300000013", 15373=>X"00000013000000130000001300000013", 15374=>X"00000013000000130000001300000013", 
15375=>X"00000013000000130000001300000013", 15376=>X"00000013000000130000001300000013", 15377=>X"00000013000000130000001300000013", 15378=>X"00000013000000130000001300000013", 15379=>X"00000013000000130000001300000013", 
15380=>X"00000013000000130000001300000013", 15381=>X"00000013000000130000001300000013", 15382=>X"00000013000000130000001300000013", 15383=>X"00000013000000130000001300000013", 15384=>X"00000013000000130000001300000013", 
15385=>X"00000013000000130000001300000013", 15386=>X"00000013000000130000001300000013", 15387=>X"00000013000000130000001300000013", 15388=>X"00000013000000130000001300000013", 15389=>X"00000013000000130000001300000013", 
15390=>X"00000013000000130000001300000013", 15391=>X"00000013000000130000001300000013", 15392=>X"00000013000000130000001300000013", 15393=>X"00000013000000130000001300000013", 15394=>X"00000013000000130000001300000013", 
15395=>X"00000013000000130000001300000013", 15396=>X"00000013000000130000001300000013", 15397=>X"00000013000000130000001300000013", 15398=>X"00000013000000130000001300000013", 15399=>X"00000013000000130000001300000013", 
15400=>X"00000013000000130000001300000013", 15401=>X"00000013000000130000001300000013", 15402=>X"00000013000000130000001300000013", 15403=>X"00000013000000130000001300000013", 15404=>X"00000013000000130000001300000013", 
15405=>X"00000013000000130000001300000013", 15406=>X"00000013000000130000001300000013", 15407=>X"00000013000000130000001300000013", 15408=>X"00000013000000130000001300000013", 15409=>X"00000013000000130000001300000013", 
15410=>X"00000013000000130000001300000013", 15411=>X"00000013000000130000001300000013", 15412=>X"00000013000000130000001300000013", 15413=>X"00000013000000130000001300000013", 15414=>X"00000013000000130000001300000013", 
15415=>X"00000013000000130000001300000013", 15416=>X"00000013000000130000001300000013", 15417=>X"00000013000000130000001300000013", 15418=>X"00000013000000130000001300000013", 15419=>X"00000013000000130000001300000013", 
15420=>X"00000013000000130000001300000013", 15421=>X"00000013000000130000001300000013", 15422=>X"00000013000000130000001300000013", 15423=>X"00000013000000130000001300000013", 15424=>X"00000013000000130000001300000013", 
15425=>X"00000013000000130000001300000013", 15426=>X"00000013000000130000001300000013", 15427=>X"00000013000000130000001300000013", 15428=>X"00000013000000130000001300000013", 15429=>X"00000013000000130000001300000013", 
15430=>X"00000013000000130000001300000013", 15431=>X"00000013000000130000001300000013", 15432=>X"00000013000000130000001300000013", 15433=>X"00000013000000130000001300000013", 15434=>X"00000013000000130000001300000013", 
15435=>X"00000013000000130000001300000013", 15436=>X"00000013000000130000001300000013", 15437=>X"00000013000000130000001300000013", 15438=>X"00000013000000130000001300000013", 15439=>X"00000013000000130000001300000013", 
15440=>X"00000013000000130000001300000013", 15441=>X"00000013000000130000001300000013", 15442=>X"00000013000000130000001300000013", 15443=>X"00000013000000130000001300000013", 15444=>X"00000013000000130000001300000013", 
15445=>X"00000013000000130000001300000013", 15446=>X"00000013000000130000001300000013", 15447=>X"00000013000000130000001300000013", 15448=>X"00000013000000130000001300000013", 15449=>X"00000013000000130000001300000013", 
15450=>X"00000013000000130000001300000013", 15451=>X"00000013000000130000001300000013", 15452=>X"00000013000000130000001300000013", 15453=>X"00000013000000130000001300000013", 15454=>X"00000013000000130000001300000013", 
15455=>X"00000013000000130000001300000013", 15456=>X"00000013000000130000001300000013", 15457=>X"00000013000000130000001300000013", 15458=>X"00000013000000130000001300000013", 15459=>X"00000013000000130000001300000013", 
15460=>X"00000013000000130000001300000013", 15461=>X"00000013000000130000001300000013", 15462=>X"00000013000000130000001300000013", 15463=>X"00000013000000130000001300000013", 15464=>X"00000013000000130000001300000013", 
15465=>X"00000013000000130000001300000013", 15466=>X"00000013000000130000001300000013", 15467=>X"00000013000000130000001300000013", 15468=>X"00000013000000130000001300000013", 15469=>X"00000013000000130000001300000013", 
15470=>X"00000013000000130000001300000013", 15471=>X"00000013000000130000001300000013", 15472=>X"00000013000000130000001300000013", 15473=>X"00000013000000130000001300000013", 15474=>X"00000013000000130000001300000013", 
15475=>X"00000013000000130000001300000013", 15476=>X"00000013000000130000001300000013", 15477=>X"00000013000000130000001300000013", 15478=>X"00000013000000130000001300000013", 15479=>X"00000013000000130000001300000013", 
15480=>X"00000013000000130000001300000013", 15481=>X"00000013000000130000001300000013", 15482=>X"00000013000000130000001300000013", 15483=>X"00000013000000130000001300000013", 15484=>X"00000013000000130000001300000013", 
15485=>X"00000013000000130000001300000013", 15486=>X"00000013000000130000001300000013", 15487=>X"00000013000000130000001300000013", 15488=>X"00000013000000130000001300000013", 15489=>X"00000013000000130000001300000013", 
15490=>X"00000013000000130000001300000013", 15491=>X"00000013000000130000001300000013", 15492=>X"00000013000000130000001300000013", 15493=>X"00000013000000130000001300000013", 15494=>X"00000013000000130000001300000013", 
15495=>X"00000013000000130000001300000013", 15496=>X"00000013000000130000001300000013", 15497=>X"00000013000000130000001300000013", 15498=>X"00000013000000130000001300000013", 15499=>X"00000013000000130000001300000013", 
15500=>X"00000013000000130000001300000013", 15501=>X"00000013000000130000001300000013", 15502=>X"00000013000000130000001300000013", 15503=>X"00000013000000130000001300000013", 15504=>X"00000013000000130000001300000013", 
15505=>X"00000013000000130000001300000013", 15506=>X"00000013000000130000001300000013", 15507=>X"00000013000000130000001300000013", 15508=>X"00000013000000130000001300000013", 15509=>X"00000013000000130000001300000013", 
15510=>X"00000013000000130000001300000013", 15511=>X"00000013000000130000001300000013", 15512=>X"00000013000000130000001300000013", 15513=>X"00000013000000130000001300000013", 15514=>X"00000013000000130000001300000013", 
15515=>X"00000013000000130000001300000013", 15516=>X"00000013000000130000001300000013", 15517=>X"00000013000000130000001300000013", 15518=>X"00000013000000130000001300000013", 15519=>X"00000013000000130000001300000013", 
15520=>X"00000013000000130000001300000013", 15521=>X"00000013000000130000001300000013", 15522=>X"00000013000000130000001300000013", 15523=>X"00000013000000130000001300000013", 15524=>X"00000013000000130000001300000013", 
15525=>X"00000013000000130000001300000013", 15526=>X"00000013000000130000001300000013", 15527=>X"00000013000000130000001300000013", 15528=>X"00000013000000130000001300000013", 15529=>X"00000013000000130000001300000013", 
15530=>X"00000013000000130000001300000013", 15531=>X"00000013000000130000001300000013", 15532=>X"00000013000000130000001300000013", 15533=>X"00000013000000130000001300000013", 15534=>X"00000013000000130000001300000013", 
15535=>X"00000013000000130000001300000013", 15536=>X"00000013000000130000001300000013", 15537=>X"00000013000000130000001300000013", 15538=>X"00000013000000130000001300000013", 15539=>X"00000013000000130000001300000013", 
15540=>X"00000013000000130000001300000013", 15541=>X"00000013000000130000001300000013", 15542=>X"00000013000000130000001300000013", 15543=>X"00000013000000130000001300000013", 15544=>X"00000013000000130000001300000013", 
15545=>X"00000013000000130000001300000013", 15546=>X"00000013000000130000001300000013", 15547=>X"00000013000000130000001300000013", 15548=>X"00000013000000130000001300000013", 15549=>X"00000013000000130000001300000013", 
15550=>X"00000013000000130000001300000013", 15551=>X"00000013000000130000001300000013", 15552=>X"00000013000000130000001300000013", 15553=>X"00000013000000130000001300000013", 15554=>X"00000013000000130000001300000013", 
15555=>X"00000013000000130000001300000013", 15556=>X"00000013000000130000001300000013", 15557=>X"00000013000000130000001300000013", 15558=>X"00000013000000130000001300000013", 15559=>X"00000013000000130000001300000013", 
15560=>X"00000013000000130000001300000013", 15561=>X"00000013000000130000001300000013", 15562=>X"00000013000000130000001300000013", 15563=>X"00000013000000130000001300000013", 15564=>X"00000013000000130000001300000013", 
15565=>X"00000013000000130000001300000013", 15566=>X"00000013000000130000001300000013", 15567=>X"00000013000000130000001300000013", 15568=>X"00000013000000130000001300000013", 15569=>X"00000013000000130000001300000013", 
15570=>X"00000013000000130000001300000013", 15571=>X"00000013000000130000001300000013", 15572=>X"00000013000000130000001300000013", 15573=>X"00000013000000130000001300000013", 15574=>X"00000013000000130000001300000013", 
15575=>X"00000013000000130000001300000013", 15576=>X"00000013000000130000001300000013", 15577=>X"00000013000000130000001300000013", 15578=>X"00000013000000130000001300000013", 15579=>X"00000013000000130000001300000013", 
15580=>X"00000013000000130000001300000013", 15581=>X"00000013000000130000001300000013", 15582=>X"00000013000000130000001300000013", 15583=>X"00000013000000130000001300000013", 15584=>X"00000013000000130000001300000013", 
15585=>X"00000013000000130000001300000013", 15586=>X"00000013000000130000001300000013", 15587=>X"00000013000000130000001300000013", 15588=>X"00000013000000130000001300000013", 15589=>X"00000013000000130000001300000013", 
15590=>X"00000013000000130000001300000013", 15591=>X"00000013000000130000001300000013", 15592=>X"00000013000000130000001300000013", 15593=>X"00000013000000130000001300000013", 15594=>X"00000013000000130000001300000013", 
15595=>X"00000013000000130000001300000013", 15596=>X"00000013000000130000001300000013", 15597=>X"00000013000000130000001300000013", 15598=>X"00000013000000130000001300000013", 15599=>X"00000013000000130000001300000013", 
15600=>X"00000013000000130000001300000013", 15601=>X"00000013000000130000001300000013", 15602=>X"00000013000000130000001300000013", 15603=>X"00000013000000130000001300000013", 15604=>X"00000013000000130000001300000013", 
15605=>X"00000013000000130000001300000013", 15606=>X"00000013000000130000001300000013", 15607=>X"00000013000000130000001300000013", 15608=>X"00000013000000130000001300000013", 15609=>X"00000013000000130000001300000013", 
15610=>X"00000013000000130000001300000013", 15611=>X"00000013000000130000001300000013", 15612=>X"00000013000000130000001300000013", 15613=>X"00000013000000130000001300000013", 15614=>X"00000013000000130000001300000013", 
15615=>X"00000013000000130000001300000013", 15616=>X"00000013000000130000001300000013", 15617=>X"00000013000000130000001300000013", 15618=>X"00000013000000130000001300000013", 15619=>X"00000013000000130000001300000013", 
15620=>X"00000013000000130000001300000013", 15621=>X"00000013000000130000001300000013", 15622=>X"00000013000000130000001300000013", 15623=>X"00000013000000130000001300000013", 15624=>X"00000013000000130000001300000013", 
15625=>X"00000013000000130000001300000013", 15626=>X"00000013000000130000001300000013", 15627=>X"00000013000000130000001300000013", 15628=>X"00000013000000130000001300000013", 15629=>X"00000013000000130000001300000013", 
15630=>X"00000013000000130000001300000013", 15631=>X"00000013000000130000001300000013", 15632=>X"00000013000000130000001300000013", 15633=>X"00000013000000130000001300000013", 15634=>X"00000013000000130000001300000013", 
15635=>X"00000013000000130000001300000013", 15636=>X"00000013000000130000001300000013", 15637=>X"00000013000000130000001300000013", 15638=>X"00000013000000130000001300000013", 15639=>X"00000013000000130000001300000013", 
15640=>X"00000013000000130000001300000013", 15641=>X"00000013000000130000001300000013", 15642=>X"00000013000000130000001300000013", 15643=>X"00000013000000130000001300000013", 15644=>X"00000013000000130000001300000013", 
15645=>X"00000013000000130000001300000013", 15646=>X"00000013000000130000001300000013", 15647=>X"00000013000000130000001300000013", 15648=>X"00000013000000130000001300000013", 15649=>X"00000013000000130000001300000013", 
15650=>X"00000013000000130000001300000013", 15651=>X"00000013000000130000001300000013", 15652=>X"00000013000000130000001300000013", 15653=>X"00000013000000130000001300000013", 15654=>X"00000013000000130000001300000013", 
15655=>X"00000013000000130000001300000013", 15656=>X"00000013000000130000001300000013", 15657=>X"00000013000000130000001300000013", 15658=>X"00000013000000130000001300000013", 15659=>X"00000013000000130000001300000013", 
15660=>X"00000013000000130000001300000013", 15661=>X"00000013000000130000001300000013", 15662=>X"00000013000000130000001300000013", 15663=>X"00000013000000130000001300000013", 15664=>X"00000013000000130000001300000013", 
15665=>X"00000013000000130000001300000013", 15666=>X"00000013000000130000001300000013", 15667=>X"00000013000000130000001300000013", 15668=>X"00000013000000130000001300000013", 15669=>X"00000013000000130000001300000013", 
15670=>X"00000013000000130000001300000013", 15671=>X"00000013000000130000001300000013", 15672=>X"00000013000000130000001300000013", 15673=>X"00000013000000130000001300000013", 15674=>X"00000013000000130000001300000013", 
15675=>X"00000013000000130000001300000013", 15676=>X"00000013000000130000001300000013", 15677=>X"00000013000000130000001300000013", 15678=>X"00000013000000130000001300000013", 15679=>X"00000013000000130000001300000013", 
15680=>X"00000013000000130000001300000013", 15681=>X"00000013000000130000001300000013", 15682=>X"00000013000000130000001300000013", 15683=>X"00000013000000130000001300000013", 15684=>X"00000013000000130000001300000013", 
15685=>X"00000013000000130000001300000013", 15686=>X"00000013000000130000001300000013", 15687=>X"00000013000000130000001300000013", 15688=>X"00000013000000130000001300000013", 15689=>X"00000013000000130000001300000013", 
15690=>X"00000013000000130000001300000013", 15691=>X"00000013000000130000001300000013", 15692=>X"00000013000000130000001300000013", 15693=>X"00000013000000130000001300000013", 15694=>X"00000013000000130000001300000013", 
15695=>X"00000013000000130000001300000013", 15696=>X"00000013000000130000001300000013", 15697=>X"00000013000000130000001300000013", 15698=>X"00000013000000130000001300000013", 15699=>X"00000013000000130000001300000013", 
15700=>X"00000013000000130000001300000013", 15701=>X"00000013000000130000001300000013", 15702=>X"00000013000000130000001300000013", 15703=>X"00000013000000130000001300000013", 15704=>X"00000013000000130000001300000013", 
15705=>X"00000013000000130000001300000013", 15706=>X"00000013000000130000001300000013", 15707=>X"00000013000000130000001300000013", 15708=>X"00000013000000130000001300000013", 15709=>X"00000013000000130000001300000013", 
15710=>X"00000013000000130000001300000013", 15711=>X"00000013000000130000001300000013", 15712=>X"00000013000000130000001300000013", 15713=>X"00000013000000130000001300000013", 15714=>X"00000013000000130000001300000013", 
15715=>X"00000013000000130000001300000013", 15716=>X"00000013000000130000001300000013", 15717=>X"00000013000000130000001300000013", 15718=>X"00000013000000130000001300000013", 15719=>X"00000013000000130000001300000013", 
15720=>X"00000013000000130000001300000013", 15721=>X"00000013000000130000001300000013", 15722=>X"00000013000000130000001300000013", 15723=>X"00000013000000130000001300000013", 15724=>X"00000013000000130000001300000013", 
15725=>X"00000013000000130000001300000013", 15726=>X"00000013000000130000001300000013", 15727=>X"00000013000000130000001300000013", 15728=>X"00000013000000130000001300000013", 15729=>X"00000013000000130000001300000013", 
15730=>X"00000013000000130000001300000013", 15731=>X"00000013000000130000001300000013", 15732=>X"00000013000000130000001300000013", 15733=>X"00000013000000130000001300000013", 15734=>X"00000013000000130000001300000013", 
15735=>X"00000013000000130000001300000013", 15736=>X"00000013000000130000001300000013", 15737=>X"00000013000000130000001300000013", 15738=>X"00000013000000130000001300000013", 15739=>X"00000013000000130000001300000013", 
15740=>X"00000013000000130000001300000013", 15741=>X"00000013000000130000001300000013", 15742=>X"00000013000000130000001300000013", 15743=>X"00000013000000130000001300000013", 15744=>X"00000013000000130000001300000013", 
15745=>X"00000013000000130000001300000013", 15746=>X"00000013000000130000001300000013", 15747=>X"00000013000000130000001300000013", 15748=>X"00000013000000130000001300000013", 15749=>X"00000013000000130000001300000013", 
15750=>X"00000013000000130000001300000013", 15751=>X"00000013000000130000001300000013", 15752=>X"00000013000000130000001300000013", 15753=>X"00000013000000130000001300000013", 15754=>X"00000013000000130000001300000013", 
15755=>X"00000013000000130000001300000013", 15756=>X"00000013000000130000001300000013", 15757=>X"00000013000000130000001300000013", 15758=>X"00000013000000130000001300000013", 15759=>X"00000013000000130000001300000013", 
15760=>X"00000013000000130000001300000013", 15761=>X"00000013000000130000001300000013", 15762=>X"00000013000000130000001300000013", 15763=>X"00000013000000130000001300000013", 15764=>X"00000013000000130000001300000013", 
15765=>X"00000013000000130000001300000013", 15766=>X"00000013000000130000001300000013", 15767=>X"00000013000000130000001300000013", 15768=>X"00000013000000130000001300000013", 15769=>X"00000013000000130000001300000013", 
15770=>X"00000013000000130000001300000013", 15771=>X"00000013000000130000001300000013", 15772=>X"00000013000000130000001300000013", 15773=>X"00000013000000130000001300000013", 15774=>X"00000013000000130000001300000013", 
15775=>X"00000013000000130000001300000013", 15776=>X"00000013000000130000001300000013", 15777=>X"00000013000000130000001300000013", 15778=>X"00000013000000130000001300000013", 15779=>X"00000013000000130000001300000013", 
15780=>X"00000013000000130000001300000013", 15781=>X"00000013000000130000001300000013", 15782=>X"00000013000000130000001300000013", 15783=>X"00000013000000130000001300000013", 15784=>X"00000013000000130000001300000013", 
15785=>X"00000013000000130000001300000013", 15786=>X"00000013000000130000001300000013", 15787=>X"00000013000000130000001300000013", 15788=>X"00000013000000130000001300000013", 15789=>X"00000013000000130000001300000013", 
15790=>X"00000013000000130000001300000013", 15791=>X"00000013000000130000001300000013", 15792=>X"00000013000000130000001300000013", 15793=>X"00000013000000130000001300000013", 15794=>X"00000013000000130000001300000013", 
15795=>X"00000013000000130000001300000013", 15796=>X"00000013000000130000001300000013", 15797=>X"00000013000000130000001300000013", 15798=>X"00000013000000130000001300000013", 15799=>X"00000013000000130000001300000013", 
15800=>X"00000013000000130000001300000013", 15801=>X"00000013000000130000001300000013", 15802=>X"00000013000000130000001300000013", 15803=>X"00000013000000130000001300000013", 15804=>X"00000013000000130000001300000013", 
15805=>X"00000013000000130000001300000013", 15806=>X"00000013000000130000001300000013", 15807=>X"00000013000000130000001300000013", 15808=>X"00000013000000130000001300000013", 15809=>X"00000013000000130000001300000013", 
15810=>X"00000013000000130000001300000013", 15811=>X"00000013000000130000001300000013", 15812=>X"00000013000000130000001300000013", 15813=>X"00000013000000130000001300000013", 15814=>X"00000013000000130000001300000013", 
15815=>X"00000013000000130000001300000013", 15816=>X"00000013000000130000001300000013", 15817=>X"00000013000000130000001300000013", 15818=>X"00000013000000130000001300000013", 15819=>X"00000013000000130000001300000013", 
15820=>X"00000013000000130000001300000013", 15821=>X"00000013000000130000001300000013", 15822=>X"00000013000000130000001300000013", 15823=>X"00000013000000130000001300000013", 15824=>X"00000013000000130000001300000013", 
15825=>X"00000013000000130000001300000013", 15826=>X"00000013000000130000001300000013", 15827=>X"00000013000000130000001300000013", 15828=>X"00000013000000130000001300000013", 15829=>X"00000013000000130000001300000013", 
15830=>X"00000013000000130000001300000013", 15831=>X"00000013000000130000001300000013", 15832=>X"00000013000000130000001300000013", 15833=>X"00000013000000130000001300000013", 15834=>X"00000013000000130000001300000013", 
15835=>X"00000013000000130000001300000013", 15836=>X"00000013000000130000001300000013", 15837=>X"00000013000000130000001300000013", 15838=>X"00000013000000130000001300000013", 15839=>X"00000013000000130000001300000013", 
15840=>X"00000013000000130000001300000013", 15841=>X"00000013000000130000001300000013", 15842=>X"00000013000000130000001300000013", 15843=>X"00000013000000130000001300000013", 15844=>X"00000013000000130000001300000013", 
15845=>X"00000013000000130000001300000013", 15846=>X"00000013000000130000001300000013", 15847=>X"00000013000000130000001300000013", 15848=>X"00000013000000130000001300000013", 15849=>X"00000013000000130000001300000013", 
15850=>X"00000013000000130000001300000013", 15851=>X"00000013000000130000001300000013", 15852=>X"00000013000000130000001300000013", 15853=>X"00000013000000130000001300000013", 15854=>X"00000013000000130000001300000013", 
15855=>X"00000013000000130000001300000013", 15856=>X"00000013000000130000001300000013", 15857=>X"00000013000000130000001300000013", 15858=>X"00000013000000130000001300000013", 15859=>X"00000013000000130000001300000013", 
15860=>X"00000013000000130000001300000013", 15861=>X"00000013000000130000001300000013", 15862=>X"00000013000000130000001300000013", 15863=>X"00000013000000130000001300000013", 15864=>X"00000013000000130000001300000013", 
15865=>X"00000013000000130000001300000013", 15866=>X"00000013000000130000001300000013", 15867=>X"00000013000000130000001300000013", 15868=>X"00000013000000130000001300000013", 15869=>X"00000013000000130000001300000013", 
15870=>X"00000013000000130000001300000013", 15871=>X"00000013000000130000001300000013", 15872=>X"00000013000000130000001300000013", 15873=>X"00000013000000130000001300000013", 15874=>X"00000013000000130000001300000013", 
15875=>X"00000013000000130000001300000013", 15876=>X"00000013000000130000001300000013", 15877=>X"00000013000000130000001300000013", 15878=>X"00000013000000130000001300000013", 15879=>X"00000013000000130000001300000013", 
15880=>X"00000013000000130000001300000013", 15881=>X"00000013000000130000001300000013", 15882=>X"00000013000000130000001300000013", 15883=>X"00000013000000130000001300000013", 15884=>X"00000013000000130000001300000013", 
15885=>X"00000013000000130000001300000013", 15886=>X"00000013000000130000001300000013", 15887=>X"00000013000000130000001300000013", 15888=>X"00000013000000130000001300000013", 15889=>X"00000013000000130000001300000013", 
15890=>X"00000013000000130000001300000013", 15891=>X"00000013000000130000001300000013", 15892=>X"00000013000000130000001300000013", 15893=>X"00000013000000130000001300000013", 15894=>X"00000013000000130000001300000013", 
15895=>X"00000013000000130000001300000013", 15896=>X"00000013000000130000001300000013", 15897=>X"00000013000000130000001300000013", 15898=>X"00000013000000130000001300000013", 15899=>X"00000013000000130000001300000013", 
15900=>X"00000013000000130000001300000013", 15901=>X"00000013000000130000001300000013", 15902=>X"00000013000000130000001300000013", 15903=>X"00000013000000130000001300000013", 15904=>X"00000013000000130000001300000013", 
15905=>X"00000013000000130000001300000013", 15906=>X"00000013000000130000001300000013", 15907=>X"00000013000000130000001300000013", 15908=>X"00000013000000130000001300000013", 15909=>X"00000013000000130000001300000013", 
15910=>X"00000013000000130000001300000013", 15911=>X"00000013000000130000001300000013", 15912=>X"00000013000000130000001300000013", 15913=>X"00000013000000130000001300000013", 15914=>X"00000013000000130000001300000013", 
15915=>X"00000013000000130000001300000013", 15916=>X"00000013000000130000001300000013", 15917=>X"00000013000000130000001300000013", 15918=>X"00000013000000130000001300000013", 15919=>X"00000013000000130000001300000013", 
15920=>X"00000013000000130000001300000013", 15921=>X"00000013000000130000001300000013", 15922=>X"00000013000000130000001300000013", 15923=>X"00000013000000130000001300000013", 15924=>X"00000013000000130000001300000013", 
15925=>X"00000013000000130000001300000013", 15926=>X"00000013000000130000001300000013", 15927=>X"00000013000000130000001300000013", 15928=>X"00000013000000130000001300000013", 15929=>X"00000013000000130000001300000013", 
15930=>X"00000013000000130000001300000013", 15931=>X"00000013000000130000001300000013", 15932=>X"00000013000000130000001300000013", 15933=>X"00000013000000130000001300000013", 15934=>X"00000013000000130000001300000013", 
15935=>X"00000013000000130000001300000013", 15936=>X"00000013000000130000001300000013", 15937=>X"00000013000000130000001300000013", 15938=>X"00000013000000130000001300000013", 15939=>X"00000013000000130000001300000013", 
15940=>X"00000013000000130000001300000013", 15941=>X"00000013000000130000001300000013", 15942=>X"00000013000000130000001300000013", 15943=>X"00000013000000130000001300000013", 15944=>X"00000013000000130000001300000013", 
15945=>X"00000013000000130000001300000013", 15946=>X"00000013000000130000001300000013", 15947=>X"00000013000000130000001300000013", 15948=>X"00000013000000130000001300000013", 15949=>X"00000013000000130000001300000013", 
15950=>X"00000013000000130000001300000013", 15951=>X"00000013000000130000001300000013", 15952=>X"00000013000000130000001300000013", 15953=>X"00000013000000130000001300000013", 15954=>X"00000013000000130000001300000013", 
15955=>X"00000013000000130000001300000013", 15956=>X"00000013000000130000001300000013", 15957=>X"00000013000000130000001300000013", 15958=>X"00000013000000130000001300000013", 15959=>X"00000013000000130000001300000013", 
15960=>X"00000013000000130000001300000013", 15961=>X"00000013000000130000001300000013", 15962=>X"00000013000000130000001300000013", 15963=>X"00000013000000130000001300000013", 15964=>X"00000013000000130000001300000013", 
15965=>X"00000013000000130000001300000013", 15966=>X"00000013000000130000001300000013", 15967=>X"00000013000000130000001300000013", 15968=>X"00000013000000130000001300000013", 15969=>X"00000013000000130000001300000013", 
15970=>X"00000013000000130000001300000013", 15971=>X"00000013000000130000001300000013", 15972=>X"00000013000000130000001300000013", 15973=>X"00000013000000130000001300000013", 15974=>X"00000013000000130000001300000013", 
15975=>X"00000013000000130000001300000013", 15976=>X"00000013000000130000001300000013", 15977=>X"00000013000000130000001300000013", 15978=>X"00000013000000130000001300000013", 15979=>X"00000013000000130000001300000013", 
15980=>X"00000013000000130000001300000013", 15981=>X"00000013000000130000001300000013", 15982=>X"00000013000000130000001300000013", 15983=>X"00000013000000130000001300000013", 15984=>X"00000013000000130000001300000013", 
15985=>X"00000013000000130000001300000013", 15986=>X"00000013000000130000001300000013", 15987=>X"00000013000000130000001300000013", 15988=>X"00000013000000130000001300000013", 15989=>X"00000013000000130000001300000013", 
15990=>X"00000013000000130000001300000013", 15991=>X"00000013000000130000001300000013", 15992=>X"00000013000000130000001300000013", 15993=>X"00000013000000130000001300000013", 15994=>X"00000013000000130000001300000013", 
15995=>X"00000013000000130000001300000013", 15996=>X"00000013000000130000001300000013", 15997=>X"00000013000000130000001300000013", 15998=>X"00000013000000130000001300000013", 15999=>X"00000013000000130000001300000013", 
16000=>X"00000013000000130000001300000013", 16001=>X"00000013000000130000001300000013", 16002=>X"00000013000000130000001300000013", 16003=>X"00000013000000130000001300000013", 16004=>X"00000013000000130000001300000013", 
16005=>X"00000013000000130000001300000013", 16006=>X"00000013000000130000001300000013", 16007=>X"00000013000000130000001300000013", 16008=>X"00000013000000130000001300000013", 16009=>X"00000013000000130000001300000013", 
16010=>X"00000013000000130000001300000013", 16011=>X"00000013000000130000001300000013", 16012=>X"00000013000000130000001300000013", 16013=>X"00000013000000130000001300000013", 16014=>X"00000013000000130000001300000013", 
16015=>X"00000013000000130000001300000013", 16016=>X"00000013000000130000001300000013", 16017=>X"00000013000000130000001300000013", 16018=>X"00000013000000130000001300000013", 16019=>X"00000013000000130000001300000013", 
16020=>X"00000013000000130000001300000013", 16021=>X"00000013000000130000001300000013", 16022=>X"00000013000000130000001300000013", 16023=>X"00000013000000130000001300000013", 16024=>X"00000013000000130000001300000013", 
16025=>X"00000013000000130000001300000013", 16026=>X"00000013000000130000001300000013", 16027=>X"00000013000000130000001300000013", 16028=>X"00000013000000130000001300000013", 16029=>X"00000013000000130000001300000013", 
16030=>X"00000013000000130000001300000013", 16031=>X"00000013000000130000001300000013", 16032=>X"00000013000000130000001300000013", 16033=>X"00000013000000130000001300000013", 16034=>X"00000013000000130000001300000013", 
16035=>X"00000013000000130000001300000013", 16036=>X"00000013000000130000001300000013", 16037=>X"00000013000000130000001300000013", 16038=>X"00000013000000130000001300000013", 16039=>X"00000012000000130000001300000013", 
16040=>X"00000012000000120000001200000012", 16041=>X"00000012000000120000001200000012", 16042=>X"00000012000000120000001200000012", 16043=>X"00000012000000120000001200000012", 16044=>X"00000012000000120000001200000012", 
16045=>X"00000012000000120000001200000012", 16046=>X"00000012000000120000001200000012", 16047=>X"00000012000000120000001200000012", 16048=>X"00000012000000120000001200000012", 16049=>X"00000012000000120000001200000012", 
16050=>X"00000012000000120000001200000012", 16051=>X"00000012000000120000001200000012", 16052=>X"00000012000000120000001200000012", 16053=>X"00000012000000120000001200000012", 16054=>X"00000012000000120000001200000012", 
16055=>X"00000012000000120000001200000012", 16056=>X"00000012000000120000001200000012", 16057=>X"00000012000000120000001200000012", 16058=>X"00000012000000120000001200000012", 16059=>X"00000012000000120000001200000012", 
16060=>X"00000012000000120000001200000012", 16061=>X"00000012000000120000001200000012", 16062=>X"00000012000000120000001200000012", 16063=>X"00000012000000120000001200000012", 16064=>X"00000012000000120000001200000012", 
16065=>X"00000012000000120000001200000012", 16066=>X"00000012000000120000001200000012", 16067=>X"00000012000000120000001200000012", 16068=>X"00000012000000120000001200000012", 16069=>X"00000012000000120000001200000012", 
16070=>X"00000012000000120000001200000012", 16071=>X"00000012000000120000001200000012", 16072=>X"00000012000000120000001200000012", 16073=>X"00000012000000120000001200000012", 16074=>X"00000012000000120000001200000012", 
16075=>X"00000012000000120000001200000012", 16076=>X"00000012000000120000001200000012", 16077=>X"00000012000000120000001200000012", 16078=>X"00000012000000120000001200000012", 16079=>X"00000012000000120000001200000012", 
16080=>X"00000012000000120000001200000012", 16081=>X"00000012000000120000001200000012", 16082=>X"00000012000000120000001200000012", 16083=>X"00000012000000120000001200000012", 16084=>X"00000012000000120000001200000012", 
16085=>X"00000012000000120000001200000012", 16086=>X"00000012000000120000001200000012", 16087=>X"00000012000000120000001200000012", 16088=>X"00000012000000120000001200000012", 16089=>X"00000012000000120000001200000012", 
16090=>X"00000012000000120000001200000012", 16091=>X"00000012000000120000001200000012", 16092=>X"00000012000000120000001200000012", 16093=>X"00000012000000120000001200000012", 16094=>X"00000012000000120000001200000012", 
16095=>X"00000012000000120000001200000012", 16096=>X"00000012000000120000001200000012", 16097=>X"00000012000000120000001200000012", 16098=>X"00000012000000120000001200000012", 16099=>X"00000012000000120000001200000012", 
16100=>X"00000012000000120000001200000012", 16101=>X"00000012000000120000001200000012", 16102=>X"00000012000000120000001200000012", 16103=>X"00000012000000120000001200000012", 16104=>X"00000012000000120000001200000012", 
16105=>X"00000012000000120000001200000012", 16106=>X"00000012000000120000001200000012", 16107=>X"00000012000000120000001200000012", 16108=>X"00000012000000120000001200000012", 16109=>X"00000012000000120000001200000012", 
16110=>X"00000012000000120000001200000012", 16111=>X"00000012000000120000001200000012", 16112=>X"00000012000000120000001200000012", 16113=>X"00000012000000120000001200000012", 16114=>X"00000012000000120000001200000012", 
16115=>X"00000012000000120000001200000012", 16116=>X"00000012000000120000001200000012", 16117=>X"00000012000000120000001200000012", 16118=>X"00000012000000120000001200000012", 16119=>X"00000012000000120000001200000012", 
16120=>X"00000012000000120000001200000012", 16121=>X"00000012000000120000001200000012", 16122=>X"00000012000000120000001200000012", 16123=>X"00000012000000120000001200000012", 16124=>X"00000012000000120000001200000012", 
16125=>X"00000012000000120000001200000012", 16126=>X"00000012000000120000001200000012", 16127=>X"00000012000000120000001200000012", 16128=>X"00000012000000120000001200000012", 16129=>X"00000012000000120000001200000012", 
16130=>X"00000012000000120000001200000012", 16131=>X"00000012000000120000001200000012", 16132=>X"00000012000000120000001200000012", 16133=>X"00000012000000120000001200000012", 16134=>X"00000012000000120000001200000012", 
16135=>X"00000012000000120000001200000012", 16136=>X"00000012000000120000001200000012", 16137=>X"00000012000000120000001200000012", 16138=>X"00000012000000120000001200000012", 16139=>X"00000012000000120000001200000012", 
16140=>X"00000012000000120000001200000012", 16141=>X"00000012000000120000001200000012", 16142=>X"00000012000000120000001200000012", 16143=>X"00000012000000120000001200000012", 16144=>X"00000012000000120000001200000012", 
16145=>X"00000012000000120000001200000012", 16146=>X"00000012000000120000001200000012", 16147=>X"00000012000000120000001200000012", 16148=>X"00000012000000120000001200000012", 16149=>X"00000012000000120000001200000012", 
16150=>X"00000012000000120000001200000012", 16151=>X"00000012000000120000001200000012", 16152=>X"00000012000000120000001200000012", 16153=>X"00000012000000120000001200000012", 16154=>X"00000012000000120000001200000012", 
16155=>X"00000012000000120000001200000012", 16156=>X"00000012000000120000001200000012", 16157=>X"00000012000000120000001200000012", 16158=>X"00000012000000120000001200000012", 16159=>X"00000012000000120000001200000012", 
16160=>X"00000012000000120000001200000012", 16161=>X"00000012000000120000001200000012", 16162=>X"00000012000000120000001200000012", 16163=>X"00000012000000120000001200000012", 16164=>X"00000012000000120000001200000012", 
16165=>X"00000012000000120000001200000012", 16166=>X"00000012000000120000001200000012", 16167=>X"00000012000000120000001200000012", 16168=>X"00000012000000120000001200000012", 16169=>X"00000012000000120000001200000012", 
16170=>X"00000012000000120000001200000012", 16171=>X"00000012000000120000001200000012", 16172=>X"00000012000000120000001200000012", 16173=>X"00000012000000120000001200000012", 16174=>X"00000012000000120000001200000012", 
16175=>X"00000012000000120000001200000012", 16176=>X"00000012000000120000001200000012", 16177=>X"00000012000000120000001200000012", 16178=>X"00000012000000120000001200000012", 16179=>X"00000012000000120000001200000012", 
16180=>X"00000012000000120000001200000012", 16181=>X"00000012000000120000001200000012", 16182=>X"00000012000000120000001200000012", 16183=>X"00000012000000120000001200000012", 16184=>X"00000012000000120000001200000012", 
16185=>X"00000012000000120000001200000012", 16186=>X"00000012000000120000001200000012", 16187=>X"00000012000000120000001200000012", 16188=>X"00000012000000120000001200000012", 16189=>X"00000012000000120000001200000012", 
16190=>X"00000012000000120000001200000012", 16191=>X"00000012000000120000001200000012", 16192=>X"00000012000000120000001200000012", 16193=>X"00000012000000120000001200000012", 16194=>X"00000012000000120000001200000012", 
16195=>X"00000012000000120000001200000012", 16196=>X"00000012000000120000001200000012", 16197=>X"00000012000000120000001200000012", 16198=>X"00000012000000120000001200000012", 16199=>X"00000012000000120000001200000012", 
16200=>X"00000012000000120000001200000012", 16201=>X"00000012000000120000001200000012", 16202=>X"00000012000000120000001200000012", 16203=>X"00000012000000120000001200000012", 16204=>X"00000012000000120000001200000012", 
16205=>X"00000012000000120000001200000012", 16206=>X"00000012000000120000001200000012", 16207=>X"00000012000000120000001200000012", 16208=>X"00000012000000120000001200000012", 16209=>X"00000012000000120000001200000012", 
16210=>X"00000012000000120000001200000012", 16211=>X"00000012000000120000001200000012", 16212=>X"00000012000000120000001200000012", 16213=>X"00000012000000120000001200000012", 16214=>X"00000012000000120000001200000012", 
16215=>X"00000012000000120000001200000012", 16216=>X"00000012000000120000001200000012", 16217=>X"00000012000000120000001200000012", 16218=>X"00000012000000120000001200000012", 16219=>X"00000012000000120000001200000012", 
16220=>X"00000012000000120000001200000012", 16221=>X"00000012000000120000001200000012", 16222=>X"00000012000000120000001200000012", 16223=>X"00000012000000120000001200000012", 16224=>X"00000012000000120000001200000012", 
16225=>X"00000012000000120000001200000012", 16226=>X"00000012000000120000001200000012", 16227=>X"00000012000000120000001200000012", 16228=>X"00000012000000120000001200000012", 16229=>X"00000012000000120000001200000012", 
16230=>X"00000012000000120000001200000012", 16231=>X"00000012000000120000001200000012", 16232=>X"00000012000000120000001200000012", 16233=>X"00000012000000120000001200000012", 16234=>X"00000012000000120000001200000012", 
16235=>X"00000012000000120000001200000012", 16236=>X"00000012000000120000001200000012", 16237=>X"00000012000000120000001200000012", 16238=>X"00000012000000120000001200000012", 16239=>X"00000012000000120000001200000012", 
16240=>X"00000012000000120000001200000012", 16241=>X"00000012000000120000001200000012", 16242=>X"00000012000000120000001200000012", 16243=>X"00000012000000120000001200000012", 16244=>X"00000012000000120000001200000012", 
16245=>X"00000012000000120000001200000012", 16246=>X"00000012000000120000001200000012", 16247=>X"00000012000000120000001200000012", 16248=>X"00000012000000120000001200000012", 16249=>X"00000012000000120000001200000012", 
16250=>X"00000012000000120000001200000012", 16251=>X"00000012000000120000001200000012", 16252=>X"00000012000000120000001200000012", 16253=>X"00000012000000120000001200000012", 16254=>X"00000012000000120000001200000012", 
16255=>X"00000012000000120000001200000012", 16256=>X"00000012000000120000001200000012", 16257=>X"00000012000000120000001200000012", 16258=>X"00000012000000120000001200000012", 16259=>X"00000012000000120000001200000012", 
16260=>X"00000012000000120000001200000012", 16261=>X"00000012000000120000001200000012", 16262=>X"00000012000000120000001200000012", 16263=>X"00000012000000120000001200000012", 16264=>X"00000012000000120000001200000012", 
16265=>X"00000012000000120000001200000012", 16266=>X"00000012000000120000001200000012", 16267=>X"00000012000000120000001200000012", 16268=>X"00000012000000120000001200000012", 16269=>X"00000012000000120000001200000012", 
16270=>X"00000012000000120000001200000012", 16271=>X"00000012000000120000001200000012", 16272=>X"00000012000000120000001200000012", 16273=>X"00000012000000120000001200000012", 16274=>X"00000012000000120000001200000012", 
16275=>X"00000012000000120000001200000012", 16276=>X"00000012000000120000001200000012", 16277=>X"00000012000000120000001200000012", 16278=>X"00000012000000120000001200000012", 16279=>X"00000012000000120000001200000012", 
16280=>X"00000012000000120000001200000012", 16281=>X"00000012000000120000001200000012", 16282=>X"00000012000000120000001200000012", 16283=>X"00000012000000120000001200000012", 16284=>X"00000012000000120000001200000012", 
16285=>X"00000012000000120000001200000012", 16286=>X"00000012000000120000001200000012", 16287=>X"00000012000000120000001200000012", 16288=>X"00000012000000120000001200000012", 16289=>X"00000012000000120000001200000012", 
16290=>X"00000012000000120000001200000012", 16291=>X"00000012000000120000001200000012", 16292=>X"00000012000000120000001200000012", 16293=>X"00000012000000120000001200000012", 16294=>X"00000012000000120000001200000012", 
16295=>X"00000012000000120000001200000012", 16296=>X"00000012000000120000001200000012", 16297=>X"00000012000000120000001200000012", 16298=>X"00000012000000120000001200000012", 16299=>X"00000012000000120000001200000012", 
16300=>X"00000012000000120000001200000012", 16301=>X"00000012000000120000001200000012", 16302=>X"00000012000000120000001200000012", 16303=>X"00000012000000120000001200000012", 16304=>X"00000012000000120000001200000012", 
16305=>X"00000012000000120000001200000012", 16306=>X"00000012000000120000001200000012", 16307=>X"00000012000000120000001200000012", 16308=>X"00000012000000120000001200000012", 16309=>X"00000012000000120000001200000012", 
16310=>X"00000012000000120000001200000012", 16311=>X"00000012000000120000001200000012", 16312=>X"00000012000000120000001200000012", 16313=>X"00000012000000120000001200000012", 16314=>X"00000012000000120000001200000012", 
16315=>X"00000012000000120000001200000012", 16316=>X"00000012000000120000001200000012", 16317=>X"00000012000000120000001200000012", 16318=>X"00000012000000120000001200000012", 16319=>X"00000012000000120000001200000012", 
16320=>X"00000012000000120000001200000012", 16321=>X"00000012000000120000001200000012", 16322=>X"00000012000000120000001200000012", 16323=>X"00000012000000120000001200000012", 16324=>X"00000012000000120000001200000012", 
16325=>X"00000012000000120000001200000012", 16326=>X"00000012000000120000001200000012", 16327=>X"00000012000000120000001200000012", 16328=>X"00000012000000120000001200000012", 16329=>X"00000012000000120000001200000012", 
16330=>X"00000012000000120000001200000012", 16331=>X"00000012000000120000001200000012", 16332=>X"00000012000000120000001200000012", 16333=>X"00000012000000120000001200000012", 16334=>X"00000012000000120000001200000012", 
16335=>X"00000012000000120000001200000012", 16336=>X"00000012000000120000001200000012", 16337=>X"00000012000000120000001200000012", 16338=>X"00000012000000120000001200000012", 16339=>X"00000012000000120000001200000012", 
16340=>X"00000012000000120000001200000012", 16341=>X"00000012000000120000001200000012", 16342=>X"00000012000000120000001200000012", 16343=>X"00000012000000120000001200000012", 16344=>X"00000012000000120000001200000012", 
16345=>X"00000012000000120000001200000012", 16346=>X"00000012000000120000001200000012", 16347=>X"00000012000000120000001200000012", 16348=>X"00000012000000120000001200000012", 16349=>X"00000012000000120000001200000012", 
16350=>X"00000012000000120000001200000012", 16351=>X"00000012000000120000001200000012", 16352=>X"00000012000000120000001200000012", 16353=>X"00000012000000120000001200000012", 16354=>X"00000012000000120000001200000012", 
16355=>X"00000012000000120000001200000012", 16356=>X"00000012000000120000001200000012", 16357=>X"00000012000000120000001200000012", 16358=>X"00000012000000120000001200000012", 16359=>X"00000012000000120000001200000012", 
16360=>X"00000012000000120000001200000012", 16361=>X"00000012000000120000001200000012", 16362=>X"00000012000000120000001200000012", 16363=>X"00000012000000120000001200000012", 16364=>X"00000012000000120000001200000012", 
16365=>X"00000012000000120000001200000012", 16366=>X"00000012000000120000001200000012", 16367=>X"00000012000000120000001200000012", 16368=>X"00000012000000120000001200000012", 16369=>X"00000012000000120000001200000012", 
16370=>X"00000012000000120000001200000012", 16371=>X"00000012000000120000001200000012", 16372=>X"00000012000000120000001200000012", 16373=>X"00000012000000120000001200000012", 16374=>X"00000012000000120000001200000012", 
16375=>X"00000012000000120000001200000012", 16376=>X"00000012000000120000001200000012", 16377=>X"00000012000000120000001200000012", 16378=>X"00000012000000120000001200000012", 16379=>X"00000012000000120000001200000012", 
16380=>X"00000012000000120000001200000012", 16381=>X"00000012000000120000001200000012", 16382=>X"00000012000000120000001200000012", 16383=>X"00000012000000120000001200000012", 16384=>X"00000012000000120000001200000012", 
16385=>X"00000012000000120000001200000012", 16386=>X"00000012000000120000001200000012", 16387=>X"00000012000000120000001200000012", 16388=>X"00000012000000120000001200000012", 16389=>X"00000012000000120000001200000012", 
16390=>X"00000012000000120000001200000012", 16391=>X"00000012000000120000001200000012", 16392=>X"00000012000000120000001200000012", 16393=>X"00000012000000120000001200000012", 16394=>X"00000012000000120000001200000012", 
16395=>X"00000012000000120000001200000012", 16396=>X"00000012000000120000001200000012", 16397=>X"00000012000000120000001200000012", 16398=>X"00000012000000120000001200000012", 16399=>X"00000012000000120000001200000012", 
16400=>X"00000012000000120000001200000012", 16401=>X"00000012000000120000001200000012", 16402=>X"00000012000000120000001200000012", 16403=>X"00000012000000120000001200000012", 16404=>X"00000012000000120000001200000012", 
16405=>X"00000012000000120000001200000012", 16406=>X"00000012000000120000001200000012", 16407=>X"00000012000000120000001200000012", 16408=>X"00000012000000120000001200000012", 16409=>X"00000012000000120000001200000012", 
16410=>X"00000012000000120000001200000012", 16411=>X"00000012000000120000001200000012", 16412=>X"00000012000000120000001200000012", 16413=>X"00000012000000120000001200000012", 16414=>X"00000012000000120000001200000012", 
16415=>X"00000012000000120000001200000012", 16416=>X"00000012000000120000001200000012", 16417=>X"00000012000000120000001200000012", 16418=>X"00000012000000120000001200000012", 16419=>X"00000012000000120000001200000012", 
16420=>X"00000012000000120000001200000012", 16421=>X"00000012000000120000001200000012", 16422=>X"00000012000000120000001200000012", 16423=>X"00000012000000120000001200000012", 16424=>X"00000012000000120000001200000012", 
16425=>X"00000012000000120000001200000012", 16426=>X"00000012000000120000001200000012", 16427=>X"00000012000000120000001200000012", 16428=>X"00000012000000120000001200000012", 16429=>X"00000012000000120000001200000012", 
16430=>X"00000012000000120000001200000012", 16431=>X"00000012000000120000001200000012", 16432=>X"00000012000000120000001200000012", 16433=>X"00000012000000120000001200000012", 16434=>X"00000012000000120000001200000012", 
16435=>X"00000012000000120000001200000012", 16436=>X"00000012000000120000001200000012", 16437=>X"00000012000000120000001200000012", 16438=>X"00000012000000120000001200000012", 16439=>X"00000012000000120000001200000012", 
16440=>X"00000012000000120000001200000012", 16441=>X"00000012000000120000001200000012", 16442=>X"00000012000000120000001200000012", 16443=>X"00000012000000120000001200000012", 16444=>X"00000012000000120000001200000012", 
16445=>X"00000012000000120000001200000012", 16446=>X"00000012000000120000001200000012", 16447=>X"00000012000000120000001200000012", 16448=>X"00000012000000120000001200000012", 16449=>X"00000012000000120000001200000012", 
16450=>X"00000012000000120000001200000012", 16451=>X"00000012000000120000001200000012", 16452=>X"00000012000000120000001200000012", 16453=>X"00000012000000120000001200000012", 16454=>X"00000012000000120000001200000012", 
16455=>X"00000012000000120000001200000012", 16456=>X"00000012000000120000001200000012", 16457=>X"00000012000000120000001200000012", 16458=>X"00000012000000120000001200000012", 16459=>X"00000012000000120000001200000012", 
16460=>X"00000012000000120000001200000012", 16461=>X"00000012000000120000001200000012", 16462=>X"00000012000000120000001200000012", 16463=>X"00000012000000120000001200000012", 16464=>X"00000012000000120000001200000012", 
16465=>X"00000012000000120000001200000012", 16466=>X"00000012000000120000001200000012", 16467=>X"00000012000000120000001200000012", 16468=>X"00000012000000120000001200000012", 16469=>X"00000012000000120000001200000012", 
16470=>X"00000012000000120000001200000012", 16471=>X"00000012000000120000001200000012", 16472=>X"00000012000000120000001200000012", 16473=>X"00000012000000120000001200000012", 16474=>X"00000012000000120000001200000012", 
16475=>X"00000012000000120000001200000012", 16476=>X"00000012000000120000001200000012", 16477=>X"00000012000000120000001200000012", 16478=>X"00000012000000120000001200000012", 16479=>X"00000012000000120000001200000012", 
16480=>X"00000012000000120000001200000012", 16481=>X"00000012000000120000001200000012", 16482=>X"00000012000000120000001200000012", 16483=>X"00000012000000120000001200000012", 16484=>X"00000012000000120000001200000012", 
16485=>X"00000012000000120000001200000012", 16486=>X"00000012000000120000001200000012", 16487=>X"00000012000000120000001200000012", 16488=>X"00000012000000120000001200000012", 16489=>X"00000012000000120000001200000012", 
16490=>X"00000012000000120000001200000012", 16491=>X"00000012000000120000001200000012", 16492=>X"00000012000000120000001200000012", 16493=>X"00000012000000120000001200000012", 16494=>X"00000012000000120000001200000012", 
16495=>X"00000012000000120000001200000012", 16496=>X"00000012000000120000001200000012", 16497=>X"00000012000000120000001200000012", 16498=>X"00000012000000120000001200000012", 16499=>X"00000012000000120000001200000012", 
16500=>X"00000012000000120000001200000012", 16501=>X"00000012000000120000001200000012", 16502=>X"00000012000000120000001200000012", 16503=>X"00000012000000120000001200000012", 16504=>X"00000012000000120000001200000012", 
16505=>X"00000012000000120000001200000012", 16506=>X"00000012000000120000001200000012", 16507=>X"00000012000000120000001200000012", 16508=>X"00000012000000120000001200000012", 16509=>X"00000012000000120000001200000012", 
16510=>X"00000012000000120000001200000012", 16511=>X"00000012000000120000001200000012", 16512=>X"00000012000000120000001200000012", 16513=>X"00000012000000120000001200000012", 16514=>X"00000012000000120000001200000012", 
16515=>X"00000012000000120000001200000012", 16516=>X"00000012000000120000001200000012", 16517=>X"00000012000000120000001200000012", 16518=>X"00000012000000120000001200000012", 16519=>X"00000012000000120000001200000012", 
16520=>X"00000012000000120000001200000012", 16521=>X"00000012000000120000001200000012", 16522=>X"00000012000000120000001200000012", 16523=>X"00000012000000120000001200000012", 16524=>X"00000012000000120000001200000012", 
16525=>X"00000012000000120000001200000012", 16526=>X"00000012000000120000001200000012", 16527=>X"00000012000000120000001200000012", 16528=>X"00000012000000120000001200000012", 16529=>X"00000012000000120000001200000012", 
16530=>X"00000012000000120000001200000012", 16531=>X"00000012000000120000001200000012", 16532=>X"00000012000000120000001200000012", 16533=>X"00000012000000120000001200000012", 16534=>X"00000012000000120000001200000012", 
16535=>X"00000012000000120000001200000012", 16536=>X"00000012000000120000001200000012", 16537=>X"00000012000000120000001200000012", 16538=>X"00000012000000120000001200000012", 16539=>X"00000012000000120000001200000012", 
16540=>X"00000012000000120000001200000012", 16541=>X"00000012000000120000001200000012", 16542=>X"00000012000000120000001200000012", 16543=>X"00000012000000120000001200000012", 16544=>X"00000012000000120000001200000012", 
16545=>X"00000012000000120000001200000012", 16546=>X"00000012000000120000001200000012", 16547=>X"00000012000000120000001200000012", 16548=>X"00000012000000120000001200000012", 16549=>X"00000012000000120000001200000012", 
16550=>X"00000012000000120000001200000012", 16551=>X"00000012000000120000001200000012", 16552=>X"00000012000000120000001200000012", 16553=>X"00000012000000120000001200000012", 16554=>X"00000012000000120000001200000012", 
16555=>X"00000012000000120000001200000012", 16556=>X"00000012000000120000001200000012", 16557=>X"00000012000000120000001200000012", 16558=>X"00000012000000120000001200000012", 16559=>X"00000012000000120000001200000012", 
16560=>X"00000012000000120000001200000012", 16561=>X"00000012000000120000001200000012", 16562=>X"00000012000000120000001200000012", 16563=>X"00000012000000120000001200000012", 16564=>X"00000012000000120000001200000012", 
16565=>X"00000012000000120000001200000012", 16566=>X"00000012000000120000001200000012", 16567=>X"00000012000000120000001200000012", 16568=>X"00000012000000120000001200000012", 16569=>X"00000012000000120000001200000012", 
16570=>X"00000012000000120000001200000012", 16571=>X"00000012000000120000001200000012", 16572=>X"00000012000000120000001200000012", 16573=>X"00000012000000120000001200000012", 16574=>X"00000012000000120000001200000012", 
16575=>X"00000012000000120000001200000012", 16576=>X"00000012000000120000001200000012", 16577=>X"00000012000000120000001200000012", 16578=>X"00000012000000120000001200000012", 16579=>X"00000012000000120000001200000012", 
16580=>X"00000012000000120000001200000012", 16581=>X"00000012000000120000001200000012", 16582=>X"00000012000000120000001200000012", 16583=>X"00000012000000120000001200000012", 16584=>X"00000012000000120000001200000012", 
16585=>X"00000012000000120000001200000012", 16586=>X"00000012000000120000001200000012", 16587=>X"00000012000000120000001200000012", 16588=>X"00000012000000120000001200000012", 16589=>X"00000012000000120000001200000012", 
16590=>X"00000012000000120000001200000012", 16591=>X"00000012000000120000001200000012", 16592=>X"00000012000000120000001200000012", 16593=>X"00000012000000120000001200000012", 16594=>X"00000012000000120000001200000012", 
16595=>X"00000012000000120000001200000012", 16596=>X"00000012000000120000001200000012", 16597=>X"00000012000000120000001200000012", 16598=>X"00000012000000120000001200000012", 16599=>X"00000012000000120000001200000012", 
16600=>X"00000012000000120000001200000012", 16601=>X"00000012000000120000001200000012", 16602=>X"00000012000000120000001200000012", 16603=>X"00000012000000120000001200000012", 16604=>X"00000012000000120000001200000012", 
16605=>X"00000012000000120000001200000012", 16606=>X"00000012000000120000001200000012", 16607=>X"00000012000000120000001200000012", 16608=>X"00000012000000120000001200000012", 16609=>X"00000012000000120000001200000012", 
16610=>X"00000012000000120000001200000012", 16611=>X"00000012000000120000001200000012", 16612=>X"00000012000000120000001200000012", 16613=>X"00000012000000120000001200000012", 16614=>X"00000012000000120000001200000012", 
16615=>X"00000012000000120000001200000012", 16616=>X"00000012000000120000001200000012", 16617=>X"00000012000000120000001200000012", 16618=>X"00000012000000120000001200000012", 16619=>X"00000012000000120000001200000012", 
16620=>X"00000012000000120000001200000012", 16621=>X"00000012000000120000001200000012", 16622=>X"00000012000000120000001200000012", 16623=>X"00000012000000120000001200000012", 16624=>X"00000012000000120000001200000012", 
16625=>X"00000012000000120000001200000012", 16626=>X"00000012000000120000001200000012", 16627=>X"00000012000000120000001200000012", 16628=>X"00000012000000120000001200000012", 16629=>X"00000012000000120000001200000012", 
16630=>X"00000012000000120000001200000012", 16631=>X"00000012000000120000001200000012", 16632=>X"00000012000000120000001200000012", 16633=>X"00000012000000120000001200000012", 16634=>X"00000012000000120000001200000012", 
16635=>X"00000012000000120000001200000012", 16636=>X"00000012000000120000001200000012", 16637=>X"00000012000000120000001200000012", 16638=>X"00000012000000120000001200000012", 16639=>X"00000012000000120000001200000012", 
16640=>X"00000012000000120000001200000012", 16641=>X"00000012000000120000001200000012", 16642=>X"00000012000000120000001200000012", 16643=>X"00000012000000120000001200000012", 16644=>X"00000012000000120000001200000012", 
16645=>X"00000012000000120000001200000012", 16646=>X"00000012000000120000001200000012", 16647=>X"00000012000000120000001200000012", 16648=>X"00000012000000120000001200000012", 16649=>X"00000012000000120000001200000012", 
16650=>X"00000012000000120000001200000012", 16651=>X"00000012000000120000001200000012", 16652=>X"00000012000000120000001200000012", 16653=>X"00000012000000120000001200000012", 16654=>X"00000012000000120000001200000012", 
16655=>X"00000012000000120000001200000012", 16656=>X"00000012000000120000001200000012", 16657=>X"00000012000000120000001200000012", 16658=>X"00000012000000120000001200000012", 16659=>X"00000012000000120000001200000012", 
16660=>X"00000012000000120000001200000012", 16661=>X"00000012000000120000001200000012", 16662=>X"00000012000000120000001200000012", 16663=>X"00000012000000120000001200000012", 16664=>X"00000012000000120000001200000012", 
16665=>X"00000012000000120000001200000012", 16666=>X"00000012000000120000001200000012", 16667=>X"00000012000000120000001200000012", 16668=>X"00000012000000120000001200000012", 16669=>X"00000012000000120000001200000012", 
16670=>X"00000012000000120000001200000012", 16671=>X"00000012000000120000001200000012", 16672=>X"00000012000000120000001200000012", 16673=>X"00000012000000120000001200000012", 16674=>X"00000012000000120000001200000012", 
16675=>X"00000012000000120000001200000012", 16676=>X"00000012000000120000001200000012", 16677=>X"00000012000000120000001200000012", 16678=>X"00000012000000120000001200000012", 16679=>X"00000012000000120000001200000012", 
16680=>X"00000012000000120000001200000012", 16681=>X"00000012000000120000001200000012", 16682=>X"00000012000000120000001200000012", 16683=>X"00000012000000120000001200000012", 16684=>X"00000012000000120000001200000012", 
16685=>X"00000012000000120000001200000012", 16686=>X"00000012000000120000001200000012", 16687=>X"00000012000000120000001200000012", 16688=>X"00000012000000120000001200000012", 16689=>X"00000012000000120000001200000012", 
16690=>X"00000012000000120000001200000012", 16691=>X"00000012000000120000001200000012", 16692=>X"00000012000000120000001200000012", 16693=>X"00000012000000120000001200000012", 16694=>X"00000012000000120000001200000012", 
16695=>X"00000012000000120000001200000012", 16696=>X"00000012000000120000001200000012", 16697=>X"00000012000000120000001200000012", 16698=>X"00000012000000120000001200000012", 16699=>X"00000012000000120000001200000012", 
16700=>X"00000012000000120000001200000012", 16701=>X"00000012000000120000001200000012", 16702=>X"00000012000000120000001200000012", 16703=>X"00000012000000120000001200000012", 16704=>X"00000012000000120000001200000012", 
16705=>X"00000012000000120000001200000012", 16706=>X"00000012000000120000001200000012", 16707=>X"00000012000000120000001200000012", 16708=>X"00000012000000120000001200000012", 16709=>X"00000012000000120000001200000012", 
16710=>X"00000012000000120000001200000012", 16711=>X"00000012000000120000001200000012", 16712=>X"00000012000000120000001200000012", 16713=>X"00000012000000120000001200000012", 16714=>X"00000012000000120000001200000012", 
16715=>X"00000012000000120000001200000012", 16716=>X"00000012000000120000001200000012", 16717=>X"00000012000000120000001200000012", 16718=>X"00000012000000120000001200000012", 16719=>X"00000012000000120000001200000012", 
16720=>X"00000012000000120000001200000012", 16721=>X"00000012000000120000001200000012", 16722=>X"00000012000000120000001200000012", 16723=>X"00000012000000120000001200000012", 16724=>X"00000012000000120000001200000012", 
16725=>X"00000012000000120000001200000012", 16726=>X"00000012000000120000001200000012", 16727=>X"00000012000000120000001200000012", 16728=>X"00000012000000120000001200000012", 16729=>X"00000012000000120000001200000012", 
16730=>X"00000012000000120000001200000012", 16731=>X"00000012000000120000001200000012", 16732=>X"00000012000000120000001200000012", 16733=>X"00000012000000120000001200000012", 16734=>X"00000012000000120000001200000012", 
16735=>X"00000012000000120000001200000012", 16736=>X"00000012000000120000001200000012", 16737=>X"00000012000000120000001200000012", 16738=>X"00000012000000120000001200000012", 16739=>X"00000012000000120000001200000012", 
16740=>X"00000012000000120000001200000012", 16741=>X"00000012000000120000001200000012", 16742=>X"00000012000000120000001200000012", 16743=>X"00000012000000120000001200000012", 16744=>X"00000012000000120000001200000012", 
16745=>X"00000012000000120000001200000012", 16746=>X"00000012000000120000001200000012", 16747=>X"00000012000000120000001200000012", 16748=>X"00000012000000120000001200000012", 16749=>X"00000012000000120000001200000012", 
16750=>X"00000012000000120000001200000012", 16751=>X"00000012000000120000001200000012", 16752=>X"00000012000000120000001200000012", 16753=>X"00000012000000120000001200000012", 16754=>X"00000012000000120000001200000012", 
16755=>X"00000012000000120000001200000012", 16756=>X"00000012000000120000001200000012", 16757=>X"00000012000000120000001200000012", 16758=>X"00000012000000120000001200000012", 16759=>X"00000012000000120000001200000012", 
16760=>X"00000012000000120000001200000012", 16761=>X"00000012000000120000001200000012", 16762=>X"00000012000000120000001200000012", 16763=>X"00000012000000120000001200000012", 16764=>X"00000012000000120000001200000012", 
16765=>X"00000012000000120000001200000012", 16766=>X"00000012000000120000001200000012", 16767=>X"00000012000000120000001200000012", 16768=>X"00000012000000120000001200000012", 16769=>X"00000012000000120000001200000012", 
16770=>X"00000012000000120000001200000012", 16771=>X"00000012000000120000001200000012", 16772=>X"00000012000000120000001200000012", 16773=>X"00000012000000120000001200000012", 16774=>X"00000012000000120000001200000012", 
16775=>X"00000012000000120000001200000012", 16776=>X"00000012000000120000001200000012", 16777=>X"00000012000000120000001200000012", 16778=>X"00000012000000120000001200000012", 16779=>X"00000012000000120000001200000012", 
16780=>X"00000012000000120000001200000012", 16781=>X"00000012000000120000001200000012", 16782=>X"00000012000000120000001200000012", 16783=>X"00000012000000120000001200000012", 16784=>X"00000012000000120000001200000012", 
16785=>X"00000012000000120000001200000012", 16786=>X"00000012000000120000001200000012", 16787=>X"00000012000000120000001200000012", 16788=>X"00000012000000120000001200000012", 16789=>X"00000012000000120000001200000012", 
16790=>X"00000012000000120000001200000012", 16791=>X"00000012000000120000001200000012", 16792=>X"00000012000000120000001200000012", 16793=>X"00000012000000120000001200000012", 16794=>X"00000012000000120000001200000012", 
16795=>X"00000012000000120000001200000012", 16796=>X"00000012000000120000001200000012", 16797=>X"00000012000000120000001200000012", 16798=>X"00000012000000120000001200000012", 16799=>X"00000012000000120000001200000012", 
16800=>X"00000012000000120000001200000012", 16801=>X"00000012000000120000001200000012", 16802=>X"00000012000000120000001200000012", 16803=>X"00000012000000120000001200000012", 16804=>X"00000012000000120000001200000012", 
16805=>X"00000012000000120000001200000012", 16806=>X"00000012000000120000001200000012", 16807=>X"00000012000000120000001200000012", 16808=>X"00000012000000120000001200000012", 16809=>X"00000012000000120000001200000012", 
16810=>X"00000012000000120000001200000012", 16811=>X"00000012000000120000001200000012", 16812=>X"00000012000000120000001200000012", 16813=>X"00000012000000120000001200000012", 16814=>X"00000012000000120000001200000012", 
16815=>X"00000012000000120000001200000012", 16816=>X"00000012000000120000001200000012", 16817=>X"00000012000000120000001200000012", 16818=>X"00000012000000120000001200000012", 16819=>X"00000012000000120000001200000012", 
16820=>X"00000012000000120000001200000012", 16821=>X"00000012000000120000001200000012", 16822=>X"00000012000000120000001200000012", 16823=>X"00000012000000120000001200000012", 16824=>X"00000012000000120000001200000012", 
16825=>X"00000012000000120000001200000012", 16826=>X"00000012000000120000001200000012", 16827=>X"00000012000000120000001200000012", 16828=>X"00000012000000120000001200000012", 16829=>X"00000012000000120000001200000012", 
16830=>X"00000012000000120000001200000012", 16831=>X"00000012000000120000001200000012", 16832=>X"00000012000000120000001200000012", 16833=>X"00000012000000120000001200000012", 16834=>X"00000012000000120000001200000012", 
16835=>X"00000012000000120000001200000012", 16836=>X"00000012000000120000001200000012", 16837=>X"00000012000000120000001200000012", 16838=>X"00000012000000120000001200000012", 16839=>X"00000012000000120000001200000012", 
16840=>X"00000012000000120000001200000012", 16841=>X"00000012000000120000001200000012", 16842=>X"00000012000000120000001200000012", 16843=>X"00000012000000120000001200000012", 16844=>X"00000012000000120000001200000012", 
16845=>X"00000012000000120000001200000012", 16846=>X"00000012000000120000001200000012", 16847=>X"00000012000000120000001200000012", 16848=>X"00000012000000120000001200000012", 16849=>X"00000011000000110000001200000012", 
16850=>X"00000011000000110000001100000011", 16851=>X"00000011000000110000001100000011", 16852=>X"00000011000000110000001100000011", 16853=>X"00000011000000110000001100000011", 16854=>X"00000011000000110000001100000011", 
16855=>X"00000011000000110000001100000011", 16856=>X"00000011000000110000001100000011", 16857=>X"00000011000000110000001100000011", 16858=>X"00000011000000110000001100000011", 16859=>X"00000011000000110000001100000011", 
16860=>X"00000011000000110000001100000011", 16861=>X"00000011000000110000001100000011", 16862=>X"00000011000000110000001100000011", 16863=>X"00000011000000110000001100000011", 16864=>X"00000011000000110000001100000011", 
16865=>X"00000011000000110000001100000011", 16866=>X"00000011000000110000001100000011", 16867=>X"00000011000000110000001100000011", 16868=>X"00000011000000110000001100000011", 16869=>X"00000011000000110000001100000011", 
16870=>X"00000011000000110000001100000011", 16871=>X"00000011000000110000001100000011", 16872=>X"00000011000000110000001100000011", 16873=>X"00000011000000110000001100000011", 16874=>X"00000011000000110000001100000011", 
16875=>X"00000011000000110000001100000011", 16876=>X"00000011000000110000001100000011", 16877=>X"00000011000000110000001100000011", 16878=>X"00000011000000110000001100000011", 16879=>X"00000011000000110000001100000011", 
16880=>X"00000011000000110000001100000011", 16881=>X"00000011000000110000001100000011", 16882=>X"00000011000000110000001100000011", 16883=>X"00000011000000110000001100000011", 16884=>X"00000011000000110000001100000011", 
16885=>X"00000011000000110000001100000011", 16886=>X"00000011000000110000001100000011", 16887=>X"00000011000000110000001100000011", 16888=>X"00000011000000110000001100000011", 16889=>X"00000011000000110000001100000011", 
16890=>X"00000011000000110000001100000011", 16891=>X"00000011000000110000001100000011", 16892=>X"00000011000000110000001100000011", 16893=>X"00000011000000110000001100000011", 16894=>X"00000011000000110000001100000011", 
16895=>X"00000011000000110000001100000011", 16896=>X"00000011000000110000001100000011", 16897=>X"00000011000000110000001100000011", 16898=>X"00000011000000110000001100000011", 16899=>X"00000011000000110000001100000011", 
16900=>X"00000011000000110000001100000011", 16901=>X"00000011000000110000001100000011", 16902=>X"00000011000000110000001100000011", 16903=>X"00000011000000110000001100000011", 16904=>X"00000011000000110000001100000011", 
16905=>X"00000011000000110000001100000011", 16906=>X"00000011000000110000001100000011", 16907=>X"00000011000000110000001100000011", 16908=>X"00000011000000110000001100000011", 16909=>X"00000011000000110000001100000011", 
16910=>X"00000011000000110000001100000011", 16911=>X"00000011000000110000001100000011", 16912=>X"00000011000000110000001100000011", 16913=>X"00000011000000110000001100000011", 16914=>X"00000011000000110000001100000011", 
16915=>X"00000011000000110000001100000011", 16916=>X"00000011000000110000001100000011", 16917=>X"00000011000000110000001100000011", 16918=>X"00000011000000110000001100000011", 16919=>X"00000011000000110000001100000011", 
16920=>X"00000011000000110000001100000011", 16921=>X"00000011000000110000001100000011", 16922=>X"00000011000000110000001100000011", 16923=>X"00000011000000110000001100000011", 16924=>X"00000011000000110000001100000011", 
16925=>X"00000011000000110000001100000011", 16926=>X"00000011000000110000001100000011", 16927=>X"00000011000000110000001100000011", 16928=>X"00000011000000110000001100000011", 16929=>X"00000011000000110000001100000011", 
16930=>X"00000011000000110000001100000011", 16931=>X"00000011000000110000001100000011", 16932=>X"00000011000000110000001100000011", 16933=>X"00000011000000110000001100000011", 16934=>X"00000011000000110000001100000011", 
16935=>X"00000011000000110000001100000011", 16936=>X"00000011000000110000001100000011", 16937=>X"00000011000000110000001100000011", 16938=>X"00000011000000110000001100000011", 16939=>X"00000011000000110000001100000011", 
16940=>X"00000011000000110000001100000011", 16941=>X"00000011000000110000001100000011", 16942=>X"00000011000000110000001100000011", 16943=>X"00000011000000110000001100000011", 16944=>X"00000011000000110000001100000011", 
16945=>X"00000011000000110000001100000011", 16946=>X"00000011000000110000001100000011", 16947=>X"00000011000000110000001100000011", 16948=>X"00000011000000110000001100000011", 16949=>X"00000011000000110000001100000011", 
16950=>X"00000011000000110000001100000011", 16951=>X"00000011000000110000001100000011", 16952=>X"00000011000000110000001100000011", 16953=>X"00000011000000110000001100000011", 16954=>X"00000011000000110000001100000011", 
16955=>X"00000011000000110000001100000011", 16956=>X"00000011000000110000001100000011", 16957=>X"00000011000000110000001100000011", 16958=>X"00000011000000110000001100000011", 16959=>X"00000011000000110000001100000011", 
16960=>X"00000011000000110000001100000011", 16961=>X"00000011000000110000001100000011", 16962=>X"00000011000000110000001100000011", 16963=>X"00000011000000110000001100000011", 16964=>X"00000011000000110000001100000011", 
16965=>X"00000011000000110000001100000011", 16966=>X"00000011000000110000001100000011", 16967=>X"00000011000000110000001100000011", 16968=>X"00000011000000110000001100000011", 16969=>X"00000011000000110000001100000011", 
16970=>X"00000011000000110000001100000011", 16971=>X"00000011000000110000001100000011", 16972=>X"00000011000000110000001100000011", 16973=>X"00000011000000110000001100000011", 16974=>X"00000011000000110000001100000011", 
16975=>X"00000011000000110000001100000011", 16976=>X"00000011000000110000001100000011", 16977=>X"00000011000000110000001100000011", 16978=>X"00000011000000110000001100000011", 16979=>X"00000011000000110000001100000011", 
16980=>X"00000011000000110000001100000011", 16981=>X"00000011000000110000001100000011", 16982=>X"00000011000000110000001100000011", 16983=>X"00000011000000110000001100000011", 16984=>X"00000011000000110000001100000011", 
16985=>X"00000011000000110000001100000011", 16986=>X"00000011000000110000001100000011", 16987=>X"00000011000000110000001100000011", 16988=>X"00000011000000110000001100000011", 16989=>X"00000011000000110000001100000011", 
16990=>X"00000011000000110000001100000011", 16991=>X"00000011000000110000001100000011", 16992=>X"00000011000000110000001100000011", 16993=>X"00000011000000110000001100000011", 16994=>X"00000011000000110000001100000011", 
16995=>X"00000011000000110000001100000011", 16996=>X"00000011000000110000001100000011", 16997=>X"00000011000000110000001100000011", 16998=>X"00000011000000110000001100000011", 16999=>X"00000011000000110000001100000011", 
17000=>X"00000011000000110000001100000011", 17001=>X"00000011000000110000001100000011", 17002=>X"00000011000000110000001100000011", 17003=>X"00000011000000110000001100000011", 17004=>X"00000011000000110000001100000011", 
17005=>X"00000011000000110000001100000011", 17006=>X"00000011000000110000001100000011", 17007=>X"00000011000000110000001100000011", 17008=>X"00000011000000110000001100000011", 17009=>X"00000011000000110000001100000011", 
17010=>X"00000011000000110000001100000011", 17011=>X"00000011000000110000001100000011", 17012=>X"00000011000000110000001100000011", 17013=>X"00000011000000110000001100000011", 17014=>X"00000011000000110000001100000011", 
17015=>X"00000011000000110000001100000011", 17016=>X"00000011000000110000001100000011", 17017=>X"00000011000000110000001100000011", 17018=>X"00000011000000110000001100000011", 17019=>X"00000011000000110000001100000011", 
17020=>X"00000011000000110000001100000011", 17021=>X"00000011000000110000001100000011", 17022=>X"00000011000000110000001100000011", 17023=>X"00000011000000110000001100000011", 17024=>X"00000011000000110000001100000011", 
17025=>X"00000011000000110000001100000011", 17026=>X"00000011000000110000001100000011", 17027=>X"00000011000000110000001100000011", 17028=>X"00000011000000110000001100000011", 17029=>X"00000011000000110000001100000011", 
17030=>X"00000011000000110000001100000011", 17031=>X"00000011000000110000001100000011", 17032=>X"00000011000000110000001100000011", 17033=>X"00000011000000110000001100000011", 17034=>X"00000011000000110000001100000011", 
17035=>X"00000011000000110000001100000011", 17036=>X"00000011000000110000001100000011", 17037=>X"00000011000000110000001100000011", 17038=>X"00000011000000110000001100000011", 17039=>X"00000011000000110000001100000011", 
17040=>X"00000011000000110000001100000011", 17041=>X"00000011000000110000001100000011", 17042=>X"00000011000000110000001100000011", 17043=>X"00000011000000110000001100000011", 17044=>X"00000011000000110000001100000011", 
17045=>X"00000011000000110000001100000011", 17046=>X"00000011000000110000001100000011", 17047=>X"00000011000000110000001100000011", 17048=>X"00000011000000110000001100000011", 17049=>X"00000011000000110000001100000011", 
17050=>X"00000011000000110000001100000011", 17051=>X"00000011000000110000001100000011", 17052=>X"00000011000000110000001100000011", 17053=>X"00000011000000110000001100000011", 17054=>X"00000011000000110000001100000011", 
17055=>X"00000011000000110000001100000011", 17056=>X"00000011000000110000001100000011", 17057=>X"00000011000000110000001100000011", 17058=>X"00000011000000110000001100000011", 17059=>X"00000011000000110000001100000011", 
17060=>X"00000011000000110000001100000011", 17061=>X"00000011000000110000001100000011", 17062=>X"00000011000000110000001100000011", 17063=>X"00000011000000110000001100000011", 17064=>X"00000011000000110000001100000011", 
17065=>X"00000011000000110000001100000011", 17066=>X"00000011000000110000001100000011", 17067=>X"00000011000000110000001100000011", 17068=>X"00000011000000110000001100000011", 17069=>X"00000011000000110000001100000011", 
17070=>X"00000011000000110000001100000011", 17071=>X"00000011000000110000001100000011", 17072=>X"00000011000000110000001100000011", 17073=>X"00000011000000110000001100000011", 17074=>X"00000011000000110000001100000011", 
17075=>X"00000011000000110000001100000011", 17076=>X"00000011000000110000001100000011", 17077=>X"00000011000000110000001100000011", 17078=>X"00000011000000110000001100000011", 17079=>X"00000011000000110000001100000011", 
17080=>X"00000011000000110000001100000011", 17081=>X"00000011000000110000001100000011", 17082=>X"00000011000000110000001100000011", 17083=>X"00000011000000110000001100000011", 17084=>X"00000011000000110000001100000011", 
17085=>X"00000011000000110000001100000011", 17086=>X"00000011000000110000001100000011", 17087=>X"00000011000000110000001100000011", 17088=>X"00000011000000110000001100000011", 17089=>X"00000011000000110000001100000011", 
17090=>X"00000011000000110000001100000011", 17091=>X"00000011000000110000001100000011", 17092=>X"00000011000000110000001100000011", 17093=>X"00000011000000110000001100000011", 17094=>X"00000011000000110000001100000011", 
17095=>X"00000011000000110000001100000011", 17096=>X"00000011000000110000001100000011", 17097=>X"00000011000000110000001100000011", 17098=>X"00000011000000110000001100000011", 17099=>X"00000011000000110000001100000011", 
17100=>X"00000011000000110000001100000011", 17101=>X"00000011000000110000001100000011", 17102=>X"00000011000000110000001100000011", 17103=>X"00000011000000110000001100000011", 17104=>X"00000011000000110000001100000011", 
17105=>X"00000011000000110000001100000011", 17106=>X"00000011000000110000001100000011", 17107=>X"00000011000000110000001100000011", 17108=>X"00000011000000110000001100000011", 17109=>X"00000011000000110000001100000011", 
17110=>X"00000011000000110000001100000011", 17111=>X"00000011000000110000001100000011", 17112=>X"00000011000000110000001100000011", 17113=>X"00000011000000110000001100000011", 17114=>X"00000011000000110000001100000011", 
17115=>X"00000011000000110000001100000011", 17116=>X"00000011000000110000001100000011", 17117=>X"00000011000000110000001100000011", 17118=>X"00000011000000110000001100000011", 17119=>X"00000011000000110000001100000011", 
17120=>X"00000011000000110000001100000011", 17121=>X"00000011000000110000001100000011", 17122=>X"00000011000000110000001100000011", 17123=>X"00000011000000110000001100000011", 17124=>X"00000011000000110000001100000011", 
17125=>X"00000011000000110000001100000011", 17126=>X"00000011000000110000001100000011", 17127=>X"00000011000000110000001100000011", 17128=>X"00000011000000110000001100000011", 17129=>X"00000011000000110000001100000011", 
17130=>X"00000011000000110000001100000011", 17131=>X"00000011000000110000001100000011", 17132=>X"00000011000000110000001100000011", 17133=>X"00000011000000110000001100000011", 17134=>X"00000011000000110000001100000011", 
17135=>X"00000011000000110000001100000011", 17136=>X"00000011000000110000001100000011", 17137=>X"00000011000000110000001100000011", 17138=>X"00000011000000110000001100000011", 17139=>X"00000011000000110000001100000011", 
17140=>X"00000011000000110000001100000011", 17141=>X"00000011000000110000001100000011", 17142=>X"00000011000000110000001100000011", 17143=>X"00000011000000110000001100000011", 17144=>X"00000011000000110000001100000011", 
17145=>X"00000011000000110000001100000011", 17146=>X"00000011000000110000001100000011", 17147=>X"00000011000000110000001100000011", 17148=>X"00000011000000110000001100000011", 17149=>X"00000011000000110000001100000011", 
17150=>X"00000011000000110000001100000011", 17151=>X"00000011000000110000001100000011", 17152=>X"00000011000000110000001100000011", 17153=>X"00000011000000110000001100000011", 17154=>X"00000011000000110000001100000011", 
17155=>X"00000011000000110000001100000011", 17156=>X"00000011000000110000001100000011", 17157=>X"00000011000000110000001100000011", 17158=>X"00000011000000110000001100000011", 17159=>X"00000011000000110000001100000011", 
17160=>X"00000011000000110000001100000011", 17161=>X"00000011000000110000001100000011", 17162=>X"00000011000000110000001100000011", 17163=>X"00000011000000110000001100000011", 17164=>X"00000011000000110000001100000011", 
17165=>X"00000011000000110000001100000011", 17166=>X"00000011000000110000001100000011", 17167=>X"00000011000000110000001100000011", 17168=>X"00000011000000110000001100000011", 17169=>X"00000011000000110000001100000011", 
17170=>X"00000011000000110000001100000011", 17171=>X"00000011000000110000001100000011", 17172=>X"00000011000000110000001100000011", 17173=>X"00000011000000110000001100000011", 17174=>X"00000011000000110000001100000011", 
17175=>X"00000011000000110000001100000011", 17176=>X"00000011000000110000001100000011", 17177=>X"00000011000000110000001100000011", 17178=>X"00000011000000110000001100000011", 17179=>X"00000011000000110000001100000011", 
17180=>X"00000011000000110000001100000011", 17181=>X"00000011000000110000001100000011", 17182=>X"00000011000000110000001100000011", 17183=>X"00000011000000110000001100000011", 17184=>X"00000011000000110000001100000011", 
17185=>X"00000011000000110000001100000011", 17186=>X"00000011000000110000001100000011", 17187=>X"00000011000000110000001100000011", 17188=>X"00000011000000110000001100000011", 17189=>X"00000011000000110000001100000011", 
17190=>X"00000011000000110000001100000011", 17191=>X"00000011000000110000001100000011", 17192=>X"00000011000000110000001100000011", 17193=>X"00000011000000110000001100000011", 17194=>X"00000011000000110000001100000011", 
17195=>X"00000011000000110000001100000011", 17196=>X"00000011000000110000001100000011", 17197=>X"00000011000000110000001100000011", 17198=>X"00000011000000110000001100000011", 17199=>X"00000011000000110000001100000011", 
17200=>X"00000011000000110000001100000011", 17201=>X"00000011000000110000001100000011", 17202=>X"00000011000000110000001100000011", 17203=>X"00000011000000110000001100000011", 17204=>X"00000011000000110000001100000011", 
17205=>X"00000011000000110000001100000011", 17206=>X"00000011000000110000001100000011", 17207=>X"00000011000000110000001100000011", 17208=>X"00000011000000110000001100000011", 17209=>X"00000011000000110000001100000011", 
17210=>X"00000011000000110000001100000011", 17211=>X"00000011000000110000001100000011", 17212=>X"00000011000000110000001100000011", 17213=>X"00000011000000110000001100000011", 17214=>X"00000011000000110000001100000011", 
17215=>X"00000011000000110000001100000011", 17216=>X"00000011000000110000001100000011", 17217=>X"00000011000000110000001100000011", 17218=>X"00000011000000110000001100000011", 17219=>X"00000011000000110000001100000011", 
17220=>X"00000011000000110000001100000011", 17221=>X"00000011000000110000001100000011", 17222=>X"00000011000000110000001100000011", 17223=>X"00000011000000110000001100000011", 17224=>X"00000011000000110000001100000011", 
17225=>X"00000011000000110000001100000011", 17226=>X"00000011000000110000001100000011", 17227=>X"00000011000000110000001100000011", 17228=>X"00000011000000110000001100000011", 17229=>X"00000011000000110000001100000011", 
17230=>X"00000011000000110000001100000011", 17231=>X"00000011000000110000001100000011", 17232=>X"00000011000000110000001100000011", 17233=>X"00000011000000110000001100000011", 17234=>X"00000011000000110000001100000011", 
17235=>X"00000011000000110000001100000011", 17236=>X"00000011000000110000001100000011", 17237=>X"00000011000000110000001100000011", 17238=>X"00000011000000110000001100000011", 17239=>X"00000011000000110000001100000011", 
17240=>X"00000011000000110000001100000011", 17241=>X"00000011000000110000001100000011", 17242=>X"00000011000000110000001100000011", 17243=>X"00000011000000110000001100000011", 17244=>X"00000011000000110000001100000011", 
17245=>X"00000011000000110000001100000011", 17246=>X"00000011000000110000001100000011", 17247=>X"00000011000000110000001100000011", 17248=>X"00000011000000110000001100000011", 17249=>X"00000011000000110000001100000011", 
17250=>X"00000011000000110000001100000011", 17251=>X"00000011000000110000001100000011", 17252=>X"00000011000000110000001100000011", 17253=>X"00000011000000110000001100000011", 17254=>X"00000011000000110000001100000011", 
17255=>X"00000011000000110000001100000011", 17256=>X"00000011000000110000001100000011", 17257=>X"00000011000000110000001100000011", 17258=>X"00000011000000110000001100000011", 17259=>X"00000011000000110000001100000011", 
17260=>X"00000011000000110000001100000011", 17261=>X"00000011000000110000001100000011", 17262=>X"00000011000000110000001100000011", 17263=>X"00000011000000110000001100000011", 17264=>X"00000011000000110000001100000011", 
17265=>X"00000011000000110000001100000011", 17266=>X"00000011000000110000001100000011", 17267=>X"00000011000000110000001100000011", 17268=>X"00000011000000110000001100000011", 17269=>X"00000011000000110000001100000011", 
17270=>X"00000011000000110000001100000011", 17271=>X"00000011000000110000001100000011", 17272=>X"00000011000000110000001100000011", 17273=>X"00000011000000110000001100000011", 17274=>X"00000011000000110000001100000011", 
17275=>X"00000011000000110000001100000011", 17276=>X"00000011000000110000001100000011", 17277=>X"00000011000000110000001100000011", 17278=>X"00000011000000110000001100000011", 17279=>X"00000011000000110000001100000011", 
17280=>X"00000011000000110000001100000011", 17281=>X"00000011000000110000001100000011", 17282=>X"00000011000000110000001100000011", 17283=>X"00000011000000110000001100000011", 17284=>X"00000011000000110000001100000011", 
17285=>X"00000011000000110000001100000011", 17286=>X"00000011000000110000001100000011", 17287=>X"00000011000000110000001100000011", 17288=>X"00000011000000110000001100000011", 17289=>X"00000011000000110000001100000011", 
17290=>X"00000011000000110000001100000011", 17291=>X"00000011000000110000001100000011", 17292=>X"00000011000000110000001100000011", 17293=>X"00000011000000110000001100000011", 17294=>X"00000011000000110000001100000011", 
17295=>X"00000011000000110000001100000011", 17296=>X"00000011000000110000001100000011", 17297=>X"00000011000000110000001100000011", 17298=>X"00000011000000110000001100000011", 17299=>X"00000011000000110000001100000011", 
17300=>X"00000011000000110000001100000011", 17301=>X"00000011000000110000001100000011", 17302=>X"00000011000000110000001100000011", 17303=>X"00000011000000110000001100000011", 17304=>X"00000011000000110000001100000011", 
17305=>X"00000011000000110000001100000011", 17306=>X"00000011000000110000001100000011", 17307=>X"00000011000000110000001100000011", 17308=>X"00000011000000110000001100000011", 17309=>X"00000011000000110000001100000011", 
17310=>X"00000011000000110000001100000011", 17311=>X"00000011000000110000001100000011", 17312=>X"00000011000000110000001100000011", 17313=>X"00000011000000110000001100000011", 17314=>X"00000011000000110000001100000011", 
17315=>X"00000011000000110000001100000011", 17316=>X"00000011000000110000001100000011", 17317=>X"00000011000000110000001100000011", 17318=>X"00000011000000110000001100000011", 17319=>X"00000011000000110000001100000011", 
17320=>X"00000011000000110000001100000011", 17321=>X"00000011000000110000001100000011", 17322=>X"00000011000000110000001100000011", 17323=>X"00000011000000110000001100000011", 17324=>X"00000011000000110000001100000011", 
17325=>X"00000011000000110000001100000011", 17326=>X"00000011000000110000001100000011", 17327=>X"00000011000000110000001100000011", 17328=>X"00000011000000110000001100000011", 17329=>X"00000011000000110000001100000011", 
17330=>X"00000011000000110000001100000011", 17331=>X"00000011000000110000001100000011", 17332=>X"00000011000000110000001100000011", 17333=>X"00000011000000110000001100000011", 17334=>X"00000011000000110000001100000011", 
17335=>X"00000011000000110000001100000011", 17336=>X"00000011000000110000001100000011", 17337=>X"00000011000000110000001100000011", 17338=>X"00000011000000110000001100000011", 17339=>X"00000011000000110000001100000011", 
17340=>X"00000011000000110000001100000011", 17341=>X"00000011000000110000001100000011", 17342=>X"00000011000000110000001100000011", 17343=>X"00000011000000110000001100000011", 17344=>X"00000011000000110000001100000011", 
17345=>X"00000011000000110000001100000011", 17346=>X"00000011000000110000001100000011", 17347=>X"00000011000000110000001100000011", 17348=>X"00000011000000110000001100000011", 17349=>X"00000011000000110000001100000011", 
17350=>X"00000011000000110000001100000011", 17351=>X"00000011000000110000001100000011", 17352=>X"00000011000000110000001100000011", 17353=>X"00000011000000110000001100000011", 17354=>X"00000011000000110000001100000011", 
17355=>X"00000011000000110000001100000011", 17356=>X"00000011000000110000001100000011", 17357=>X"00000011000000110000001100000011", 17358=>X"00000011000000110000001100000011", 17359=>X"00000011000000110000001100000011", 
17360=>X"00000011000000110000001100000011", 17361=>X"00000011000000110000001100000011", 17362=>X"00000011000000110000001100000011", 17363=>X"00000011000000110000001100000011", 17364=>X"00000011000000110000001100000011", 
17365=>X"00000011000000110000001100000011", 17366=>X"00000011000000110000001100000011", 17367=>X"00000011000000110000001100000011", 17368=>X"00000011000000110000001100000011", 17369=>X"00000011000000110000001100000011", 
17370=>X"00000011000000110000001100000011", 17371=>X"00000011000000110000001100000011", 17372=>X"00000011000000110000001100000011", 17373=>X"00000011000000110000001100000011", 17374=>X"00000011000000110000001100000011", 
17375=>X"00000011000000110000001100000011", 17376=>X"00000011000000110000001100000011", 17377=>X"00000011000000110000001100000011", 17378=>X"00000011000000110000001100000011", 17379=>X"00000011000000110000001100000011", 
17380=>X"00000011000000110000001100000011", 17381=>X"00000011000000110000001100000011", 17382=>X"00000011000000110000001100000011", 17383=>X"00000011000000110000001100000011", 17384=>X"00000011000000110000001100000011", 
17385=>X"00000011000000110000001100000011", 17386=>X"00000011000000110000001100000011", 17387=>X"00000011000000110000001100000011", 17388=>X"00000011000000110000001100000011", 17389=>X"00000011000000110000001100000011", 
17390=>X"00000011000000110000001100000011", 17391=>X"00000011000000110000001100000011", 17392=>X"00000011000000110000001100000011", 17393=>X"00000011000000110000001100000011", 17394=>X"00000011000000110000001100000011", 
17395=>X"00000011000000110000001100000011", 17396=>X"00000011000000110000001100000011", 17397=>X"00000011000000110000001100000011", 17398=>X"00000011000000110000001100000011", 17399=>X"00000011000000110000001100000011", 
17400=>X"00000011000000110000001100000011", 17401=>X"00000011000000110000001100000011", 17402=>X"00000011000000110000001100000011", 17403=>X"00000011000000110000001100000011", 17404=>X"00000011000000110000001100000011", 
17405=>X"00000011000000110000001100000011", 17406=>X"00000011000000110000001100000011", 17407=>X"00000011000000110000001100000011", 17408=>X"00000011000000110000001100000011", 17409=>X"00000011000000110000001100000011", 
17410=>X"00000011000000110000001100000011", 17411=>X"00000011000000110000001100000011", 17412=>X"00000011000000110000001100000011", 17413=>X"00000011000000110000001100000011", 17414=>X"00000011000000110000001100000011", 
17415=>X"00000011000000110000001100000011", 17416=>X"00000011000000110000001100000011", 17417=>X"00000011000000110000001100000011", 17418=>X"00000011000000110000001100000011", 17419=>X"00000011000000110000001100000011", 
17420=>X"00000011000000110000001100000011", 17421=>X"00000011000000110000001100000011", 17422=>X"00000011000000110000001100000011", 17423=>X"00000011000000110000001100000011", 17424=>X"00000011000000110000001100000011", 
17425=>X"00000011000000110000001100000011", 17426=>X"00000011000000110000001100000011", 17427=>X"00000011000000110000001100000011", 17428=>X"00000011000000110000001100000011", 17429=>X"00000011000000110000001100000011", 
17430=>X"00000011000000110000001100000011", 17431=>X"00000011000000110000001100000011", 17432=>X"00000011000000110000001100000011", 17433=>X"00000011000000110000001100000011", 17434=>X"00000011000000110000001100000011", 
17435=>X"00000011000000110000001100000011", 17436=>X"00000011000000110000001100000011", 17437=>X"00000011000000110000001100000011", 17438=>X"00000011000000110000001100000011", 17439=>X"00000011000000110000001100000011", 
17440=>X"00000011000000110000001100000011", 17441=>X"00000011000000110000001100000011", 17442=>X"00000011000000110000001100000011", 17443=>X"00000011000000110000001100000011", 17444=>X"00000011000000110000001100000011", 
17445=>X"00000011000000110000001100000011", 17446=>X"00000011000000110000001100000011", 17447=>X"00000011000000110000001100000011", 17448=>X"00000011000000110000001100000011", 17449=>X"00000011000000110000001100000011", 
17450=>X"00000011000000110000001100000011", 17451=>X"00000011000000110000001100000011", 17452=>X"00000011000000110000001100000011", 17453=>X"00000011000000110000001100000011", 17454=>X"00000011000000110000001100000011", 
17455=>X"00000011000000110000001100000011", 17456=>X"00000011000000110000001100000011", 17457=>X"00000011000000110000001100000011", 17458=>X"00000011000000110000001100000011", 17459=>X"00000011000000110000001100000011", 
17460=>X"00000011000000110000001100000011", 17461=>X"00000011000000110000001100000011", 17462=>X"00000011000000110000001100000011", 17463=>X"00000011000000110000001100000011", 17464=>X"00000011000000110000001100000011", 
17465=>X"00000011000000110000001100000011", 17466=>X"00000011000000110000001100000011", 17467=>X"00000011000000110000001100000011", 17468=>X"00000011000000110000001100000011", 17469=>X"00000011000000110000001100000011", 
17470=>X"00000011000000110000001100000011", 17471=>X"00000011000000110000001100000011", 17472=>X"00000011000000110000001100000011", 17473=>X"00000011000000110000001100000011", 17474=>X"00000011000000110000001100000011", 
17475=>X"00000011000000110000001100000011", 17476=>X"00000011000000110000001100000011", 17477=>X"00000011000000110000001100000011", 17478=>X"00000011000000110000001100000011", 17479=>X"00000011000000110000001100000011", 
17480=>X"00000011000000110000001100000011", 17481=>X"00000011000000110000001100000011", 17482=>X"00000011000000110000001100000011", 17483=>X"00000011000000110000001100000011", 17484=>X"00000011000000110000001100000011", 
17485=>X"00000011000000110000001100000011", 17486=>X"00000011000000110000001100000011", 17487=>X"00000011000000110000001100000011", 17488=>X"00000011000000110000001100000011", 17489=>X"00000011000000110000001100000011", 
17490=>X"00000011000000110000001100000011", 17491=>X"00000011000000110000001100000011", 17492=>X"00000011000000110000001100000011", 17493=>X"00000011000000110000001100000011", 17494=>X"00000011000000110000001100000011", 
17495=>X"00000011000000110000001100000011", 17496=>X"00000011000000110000001100000011", 17497=>X"00000011000000110000001100000011", 17498=>X"00000011000000110000001100000011", 17499=>X"00000011000000110000001100000011", 
17500=>X"00000011000000110000001100000011", 17501=>X"00000011000000110000001100000011", 17502=>X"00000011000000110000001100000011", 17503=>X"00000011000000110000001100000011", 17504=>X"00000011000000110000001100000011", 
17505=>X"00000011000000110000001100000011", 17506=>X"00000011000000110000001100000011", 17507=>X"00000011000000110000001100000011", 17508=>X"00000011000000110000001100000011", 17509=>X"00000011000000110000001100000011", 
17510=>X"00000011000000110000001100000011", 17511=>X"00000011000000110000001100000011", 17512=>X"00000011000000110000001100000011", 17513=>X"00000011000000110000001100000011", 17514=>X"00000011000000110000001100000011", 
17515=>X"00000011000000110000001100000011", 17516=>X"00000011000000110000001100000011", 17517=>X"00000011000000110000001100000011", 17518=>X"00000011000000110000001100000011", 17519=>X"00000011000000110000001100000011", 
17520=>X"00000011000000110000001100000011", 17521=>X"00000011000000110000001100000011", 17522=>X"00000011000000110000001100000011", 17523=>X"00000011000000110000001100000011", 17524=>X"00000011000000110000001100000011", 
17525=>X"00000011000000110000001100000011", 17526=>X"00000011000000110000001100000011", 17527=>X"00000011000000110000001100000011", 17528=>X"00000011000000110000001100000011", 17529=>X"00000011000000110000001100000011", 
17530=>X"00000011000000110000001100000011", 17531=>X"00000011000000110000001100000011", 17532=>X"00000011000000110000001100000011", 17533=>X"00000011000000110000001100000011", 17534=>X"00000011000000110000001100000011", 
17535=>X"00000011000000110000001100000011", 17536=>X"00000011000000110000001100000011", 17537=>X"00000011000000110000001100000011", 17538=>X"00000011000000110000001100000011", 17539=>X"00000011000000110000001100000011", 
17540=>X"00000011000000110000001100000011", 17541=>X"00000011000000110000001100000011", 17542=>X"00000011000000110000001100000011", 17543=>X"00000011000000110000001100000011", 17544=>X"00000011000000110000001100000011", 
17545=>X"00000011000000110000001100000011", 17546=>X"00000011000000110000001100000011", 17547=>X"00000011000000110000001100000011", 17548=>X"00000011000000110000001100000011", 17549=>X"00000011000000110000001100000011", 
17550=>X"00000011000000110000001100000011", 17551=>X"00000011000000110000001100000011", 17552=>X"00000011000000110000001100000011", 17553=>X"00000011000000110000001100000011", 17554=>X"00000011000000110000001100000011", 
17555=>X"00000011000000110000001100000011", 17556=>X"00000011000000110000001100000011", 17557=>X"00000011000000110000001100000011", 17558=>X"00000011000000110000001100000011", 17559=>X"00000011000000110000001100000011", 
17560=>X"00000011000000110000001100000011", 17561=>X"00000011000000110000001100000011", 17562=>X"00000011000000110000001100000011", 17563=>X"00000011000000110000001100000011", 17564=>X"00000011000000110000001100000011", 
17565=>X"00000011000000110000001100000011", 17566=>X"00000011000000110000001100000011", 17567=>X"00000011000000110000001100000011", 17568=>X"00000011000000110000001100000011", 17569=>X"00000011000000110000001100000011", 
17570=>X"00000011000000110000001100000011", 17571=>X"00000011000000110000001100000011", 17572=>X"00000011000000110000001100000011", 17573=>X"00000011000000110000001100000011", 17574=>X"00000011000000110000001100000011", 
17575=>X"00000011000000110000001100000011", 17576=>X"00000011000000110000001100000011", 17577=>X"00000011000000110000001100000011", 17578=>X"00000011000000110000001100000011", 17579=>X"00000011000000110000001100000011", 
17580=>X"00000011000000110000001100000011", 17581=>X"00000011000000110000001100000011", 17582=>X"00000011000000110000001100000011", 17583=>X"00000011000000110000001100000011", 17584=>X"00000011000000110000001100000011", 
17585=>X"00000011000000110000001100000011", 17586=>X"00000011000000110000001100000011", 17587=>X"00000011000000110000001100000011", 17588=>X"00000011000000110000001100000011", 17589=>X"00000011000000110000001100000011", 
17590=>X"00000011000000110000001100000011", 17591=>X"00000011000000110000001100000011", 17592=>X"00000011000000110000001100000011", 17593=>X"00000011000000110000001100000011", 17594=>X"00000011000000110000001100000011", 
17595=>X"00000011000000110000001100000011", 17596=>X"00000011000000110000001100000011", 17597=>X"00000011000000110000001100000011", 17598=>X"00000011000000110000001100000011", 17599=>X"00000011000000110000001100000011", 
17600=>X"00000011000000110000001100000011", 17601=>X"00000011000000110000001100000011", 17602=>X"00000011000000110000001100000011", 17603=>X"00000011000000110000001100000011", 17604=>X"00000011000000110000001100000011", 
17605=>X"00000011000000110000001100000011", 17606=>X"00000011000000110000001100000011", 17607=>X"00000011000000110000001100000011", 17608=>X"00000011000000110000001100000011", 17609=>X"00000011000000110000001100000011", 
17610=>X"00000011000000110000001100000011", 17611=>X"00000011000000110000001100000011", 17612=>X"00000011000000110000001100000011", 17613=>X"00000011000000110000001100000011", 17614=>X"00000011000000110000001100000011", 
17615=>X"00000011000000110000001100000011", 17616=>X"00000011000000110000001100000011", 17617=>X"00000011000000110000001100000011", 17618=>X"00000011000000110000001100000011", 17619=>X"00000011000000110000001100000011", 
17620=>X"00000011000000110000001100000011", 17621=>X"00000011000000110000001100000011", 17622=>X"00000011000000110000001100000011", 17623=>X"00000011000000110000001100000011", 17624=>X"00000011000000110000001100000011", 
17625=>X"00000011000000110000001100000011", 17626=>X"00000011000000110000001100000011", 17627=>X"00000011000000110000001100000011", 17628=>X"00000011000000110000001100000011", 17629=>X"00000011000000110000001100000011", 
17630=>X"00000011000000110000001100000011", 17631=>X"00000011000000110000001100000011", 17632=>X"00000011000000110000001100000011", 17633=>X"00000011000000110000001100000011", 17634=>X"00000011000000110000001100000011", 
17635=>X"00000011000000110000001100000011", 17636=>X"00000011000000110000001100000011", 17637=>X"00000011000000110000001100000011", 17638=>X"00000011000000110000001100000011", 17639=>X"00000011000000110000001100000011", 
17640=>X"00000011000000110000001100000011", 17641=>X"00000011000000110000001100000011", 17642=>X"00000011000000110000001100000011", 17643=>X"00000011000000110000001100000011", 17644=>X"00000011000000110000001100000011", 
17645=>X"00000011000000110000001100000011", 17646=>X"00000011000000110000001100000011", 17647=>X"00000011000000110000001100000011", 17648=>X"00000011000000110000001100000011", 17649=>X"00000011000000110000001100000011", 
17650=>X"00000011000000110000001100000011", 17651=>X"00000011000000110000001100000011", 17652=>X"00000011000000110000001100000011", 17653=>X"00000011000000110000001100000011", 17654=>X"00000011000000110000001100000011", 
17655=>X"00000011000000110000001100000011", 17656=>X"00000011000000110000001100000011", 17657=>X"00000011000000110000001100000011", 17658=>X"00000011000000110000001100000011", 17659=>X"00000011000000110000001100000011", 
17660=>X"00000011000000110000001100000011", 17661=>X"00000011000000110000001100000011", 17662=>X"00000011000000110000001100000011", 17663=>X"00000011000000110000001100000011", 17664=>X"00000011000000110000001100000011", 
17665=>X"00000011000000110000001100000011", 17666=>X"00000011000000110000001100000011", 17667=>X"00000011000000110000001100000011", 17668=>X"00000011000000110000001100000011", 17669=>X"00000011000000110000001100000011", 
17670=>X"00000011000000110000001100000011", 17671=>X"00000011000000110000001100000011", 17672=>X"00000011000000110000001100000011", 17673=>X"00000011000000110000001100000011", 17674=>X"00000011000000110000001100000011", 
17675=>X"00000011000000110000001100000011", 17676=>X"00000011000000110000001100000011", 17677=>X"00000011000000110000001100000011", 17678=>X"00000011000000110000001100000011", 17679=>X"00000011000000110000001100000011", 
17680=>X"00000011000000110000001100000011", 17681=>X"00000011000000110000001100000011", 17682=>X"00000011000000110000001100000011", 17683=>X"00000011000000110000001100000011", 17684=>X"00000011000000110000001100000011", 
17685=>X"00000011000000110000001100000011", 17686=>X"00000011000000110000001100000011", 17687=>X"00000011000000110000001100000011", 17688=>X"00000011000000110000001100000011", 17689=>X"00000011000000110000001100000011", 
17690=>X"00000011000000110000001100000011", 17691=>X"00000011000000110000001100000011", 17692=>X"00000011000000110000001100000011", 17693=>X"00000011000000110000001100000011", 17694=>X"00000011000000110000001100000011", 
17695=>X"00000011000000110000001100000011", 17696=>X"00000011000000110000001100000011", 17697=>X"00000011000000110000001100000011", 17698=>X"00000011000000110000001100000011", 17699=>X"00000011000000110000001100000011", 
17700=>X"00000011000000110000001100000011", 17701=>X"00000011000000110000001100000011", 17702=>X"00000011000000110000001100000011", 17703=>X"00000011000000110000001100000011", 17704=>X"00000011000000110000001100000011", 
17705=>X"00000011000000110000001100000011", 17706=>X"00000011000000110000001100000011", 17707=>X"00000011000000110000001100000011", 17708=>X"00000011000000110000001100000011", 17709=>X"00000011000000110000001100000011", 
17710=>X"00000011000000110000001100000011", 17711=>X"00000011000000110000001100000011", 17712=>X"00000011000000110000001100000011", 17713=>X"00000011000000110000001100000011", 17714=>X"00000011000000110000001100000011", 
17715=>X"00000011000000110000001100000011", 17716=>X"00000011000000110000001100000011", 17717=>X"00000011000000110000001100000011", 17718=>X"00000011000000110000001100000011", 17719=>X"00000011000000110000001100000011", 
17720=>X"00000011000000110000001100000011", 17721=>X"00000011000000110000001100000011", 17722=>X"00000011000000110000001100000011", 17723=>X"00000011000000110000001100000011", 17724=>X"00000011000000110000001100000011", 
17725=>X"00000011000000110000001100000011", 17726=>X"00000011000000110000001100000011", 17727=>X"00000011000000110000001100000011", 17728=>X"00000011000000110000001100000011", 17729=>X"00000011000000110000001100000011", 
17730=>X"00000011000000110000001100000011", 17731=>X"00000011000000110000001100000011", 17732=>X"00000011000000110000001100000011", 17733=>X"00000011000000110000001100000011", 17734=>X"00000011000000110000001100000011", 
17735=>X"00000011000000110000001100000011", 17736=>X"00000011000000110000001100000011", 17737=>X"00000011000000110000001100000011", 17738=>X"00000011000000110000001100000011", 17739=>X"00000011000000110000001100000011", 
17740=>X"00000011000000110000001100000011", 17741=>X"00000011000000110000001100000011", 17742=>X"00000011000000110000001100000011", 17743=>X"00000011000000110000001100000011", 17744=>X"00000011000000110000001100000011", 
17745=>X"00000011000000110000001100000011", 17746=>X"00000011000000110000001100000011", 17747=>X"00000011000000110000001100000011", 17748=>X"00000011000000110000001100000011", 17749=>X"00000011000000110000001100000011", 
17750=>X"00000011000000110000001100000011", 17751=>X"00000011000000110000001100000011", 17752=>X"00000011000000110000001100000011", 17753=>X"00000011000000110000001100000011", 17754=>X"00000011000000110000001100000011", 
17755=>X"00000011000000110000001100000011", 17756=>X"00000011000000110000001100000011", 17757=>X"00000010000000100000001100000011", 17758=>X"00000010000000100000001000000010", 17759=>X"00000010000000100000001000000010", 
17760=>X"00000010000000100000001000000010", 17761=>X"00000010000000100000001000000010", 17762=>X"00000010000000100000001000000010", 17763=>X"00000010000000100000001000000010", 17764=>X"00000010000000100000001000000010", 
17765=>X"00000010000000100000001000000010", 17766=>X"00000010000000100000001000000010", 17767=>X"00000010000000100000001000000010", 17768=>X"00000010000000100000001000000010", 17769=>X"00000010000000100000001000000010", 
17770=>X"00000010000000100000001000000010", 17771=>X"00000010000000100000001000000010", 17772=>X"00000010000000100000001000000010", 17773=>X"00000010000000100000001000000010", 17774=>X"00000010000000100000001000000010", 
17775=>X"00000010000000100000001000000010", 17776=>X"00000010000000100000001000000010", 17777=>X"00000010000000100000001000000010", 17778=>X"00000010000000100000001000000010", 17779=>X"00000010000000100000001000000010", 
17780=>X"00000010000000100000001000000010", 17781=>X"00000010000000100000001000000010", 17782=>X"00000010000000100000001000000010", 17783=>X"00000010000000100000001000000010", 17784=>X"00000010000000100000001000000010", 
17785=>X"00000010000000100000001000000010", 17786=>X"00000010000000100000001000000010", 17787=>X"00000010000000100000001000000010", 17788=>X"00000010000000100000001000000010", 17789=>X"00000010000000100000001000000010", 
17790=>X"00000010000000100000001000000010", 17791=>X"00000010000000100000001000000010", 17792=>X"00000010000000100000001000000010", 17793=>X"00000010000000100000001000000010", 17794=>X"00000010000000100000001000000010", 
17795=>X"00000010000000100000001000000010", 17796=>X"00000010000000100000001000000010", 17797=>X"00000010000000100000001000000010", 17798=>X"00000010000000100000001000000010", 17799=>X"00000010000000100000001000000010", 
17800=>X"00000010000000100000001000000010", 17801=>X"00000010000000100000001000000010", 17802=>X"00000010000000100000001000000010", 17803=>X"00000010000000100000001000000010", 17804=>X"00000010000000100000001000000010", 
17805=>X"00000010000000100000001000000010", 17806=>X"00000010000000100000001000000010", 17807=>X"00000010000000100000001000000010", 17808=>X"00000010000000100000001000000010", 17809=>X"00000010000000100000001000000010", 
17810=>X"00000010000000100000001000000010", 17811=>X"00000010000000100000001000000010", 17812=>X"00000010000000100000001000000010", 17813=>X"00000010000000100000001000000010", 17814=>X"00000010000000100000001000000010", 
17815=>X"00000010000000100000001000000010", 17816=>X"00000010000000100000001000000010", 17817=>X"00000010000000100000001000000010", 17818=>X"00000010000000100000001000000010", 17819=>X"00000010000000100000001000000010", 
17820=>X"00000010000000100000001000000010", 17821=>X"00000010000000100000001000000010", 17822=>X"00000010000000100000001000000010", 17823=>X"00000010000000100000001000000010", 17824=>X"00000010000000100000001000000010", 
17825=>X"00000010000000100000001000000010", 17826=>X"00000010000000100000001000000010", 17827=>X"00000010000000100000001000000010", 17828=>X"00000010000000100000001000000010", 17829=>X"00000010000000100000001000000010", 
17830=>X"00000010000000100000001000000010", 17831=>X"00000010000000100000001000000010", 17832=>X"00000010000000100000001000000010", 17833=>X"00000010000000100000001000000010", 17834=>X"00000010000000100000001000000010", 
17835=>X"00000010000000100000001000000010", 17836=>X"00000010000000100000001000000010", 17837=>X"00000010000000100000001000000010", 17838=>X"00000010000000100000001000000010", 17839=>X"00000010000000100000001000000010", 
17840=>X"00000010000000100000001000000010", 17841=>X"00000010000000100000001000000010", 17842=>X"00000010000000100000001000000010", 17843=>X"00000010000000100000001000000010", 17844=>X"00000010000000100000001000000010", 
17845=>X"00000010000000100000001000000010", 17846=>X"00000010000000100000001000000010", 17847=>X"00000010000000100000001000000010", 17848=>X"00000010000000100000001000000010", 17849=>X"00000010000000100000001000000010", 
17850=>X"00000010000000100000001000000010", 17851=>X"00000010000000100000001000000010", 17852=>X"00000010000000100000001000000010", 17853=>X"00000010000000100000001000000010", 17854=>X"00000010000000100000001000000010", 
17855=>X"00000010000000100000001000000010", 17856=>X"00000010000000100000001000000010", 17857=>X"00000010000000100000001000000010", 17858=>X"00000010000000100000001000000010", 17859=>X"00000010000000100000001000000010", 
17860=>X"00000010000000100000001000000010", 17861=>X"00000010000000100000001000000010", 17862=>X"00000010000000100000001000000010", 17863=>X"00000010000000100000001000000010", 17864=>X"00000010000000100000001000000010", 
17865=>X"00000010000000100000001000000010", 17866=>X"00000010000000100000001000000010", 17867=>X"00000010000000100000001000000010", 17868=>X"00000010000000100000001000000010", 17869=>X"00000010000000100000001000000010", 
17870=>X"00000010000000100000001000000010", 17871=>X"00000010000000100000001000000010", 17872=>X"00000010000000100000001000000010", 17873=>X"00000010000000100000001000000010", 17874=>X"00000010000000100000001000000010", 
17875=>X"00000010000000100000001000000010", 17876=>X"00000010000000100000001000000010", 17877=>X"00000010000000100000001000000010", 17878=>X"00000010000000100000001000000010", 17879=>X"00000010000000100000001000000010", 
17880=>X"00000010000000100000001000000010", 17881=>X"00000010000000100000001000000010", 17882=>X"00000010000000100000001000000010", 17883=>X"00000010000000100000001000000010", 17884=>X"00000010000000100000001000000010", 
17885=>X"00000010000000100000001000000010", 17886=>X"00000010000000100000001000000010", 17887=>X"00000010000000100000001000000010", 17888=>X"00000010000000100000001000000010", 17889=>X"00000010000000100000001000000010", 
17890=>X"00000010000000100000001000000010", 17891=>X"00000010000000100000001000000010", 17892=>X"00000010000000100000001000000010", 17893=>X"00000010000000100000001000000010", 17894=>X"00000010000000100000001000000010", 
17895=>X"00000010000000100000001000000010", 17896=>X"00000010000000100000001000000010", 17897=>X"00000010000000100000001000000010", 17898=>X"00000010000000100000001000000010", 17899=>X"00000010000000100000001000000010", 
17900=>X"00000010000000100000001000000010", 17901=>X"00000010000000100000001000000010", 17902=>X"00000010000000100000001000000010", 17903=>X"00000010000000100000001000000010", 17904=>X"00000010000000100000001000000010", 
17905=>X"00000010000000100000001000000010", 17906=>X"00000010000000100000001000000010", 17907=>X"00000010000000100000001000000010", 17908=>X"00000010000000100000001000000010", 17909=>X"00000010000000100000001000000010", 
17910=>X"00000010000000100000001000000010", 17911=>X"00000010000000100000001000000010", 17912=>X"00000010000000100000001000000010", 17913=>X"00000010000000100000001000000010", 17914=>X"00000010000000100000001000000010", 
17915=>X"00000010000000100000001000000010", 17916=>X"00000010000000100000001000000010", 17917=>X"00000010000000100000001000000010", 17918=>X"00000010000000100000001000000010", 17919=>X"00000010000000100000001000000010", 
17920=>X"00000010000000100000001000000010", 17921=>X"00000010000000100000001000000010", 17922=>X"00000010000000100000001000000010", 17923=>X"00000010000000100000001000000010", 17924=>X"00000010000000100000001000000010", 
17925=>X"00000010000000100000001000000010", 17926=>X"00000010000000100000001000000010", 17927=>X"00000010000000100000001000000010", 17928=>X"00000010000000100000001000000010", 17929=>X"00000010000000100000001000000010", 
17930=>X"00000010000000100000001000000010", 17931=>X"00000010000000100000001000000010", 17932=>X"00000010000000100000001000000010", 17933=>X"00000010000000100000001000000010", 17934=>X"00000010000000100000001000000010", 
17935=>X"00000010000000100000001000000010", 17936=>X"00000010000000100000001000000010", 17937=>X"00000010000000100000001000000010", 17938=>X"00000010000000100000001000000010", 17939=>X"00000010000000100000001000000010", 
17940=>X"00000010000000100000001000000010", 17941=>X"00000010000000100000001000000010", 17942=>X"00000010000000100000001000000010", 17943=>X"00000010000000100000001000000010", 17944=>X"00000010000000100000001000000010", 
17945=>X"00000010000000100000001000000010", 17946=>X"00000010000000100000001000000010", 17947=>X"00000010000000100000001000000010", 17948=>X"00000010000000100000001000000010", 17949=>X"00000010000000100000001000000010", 
17950=>X"00000010000000100000001000000010", 17951=>X"00000010000000100000001000000010", 17952=>X"00000010000000100000001000000010", 17953=>X"00000010000000100000001000000010", 17954=>X"00000010000000100000001000000010", 
17955=>X"00000010000000100000001000000010", 17956=>X"00000010000000100000001000000010", 17957=>X"00000010000000100000001000000010", 17958=>X"00000010000000100000001000000010", 17959=>X"00000010000000100000001000000010", 
17960=>X"00000010000000100000001000000010", 17961=>X"00000010000000100000001000000010", 17962=>X"00000010000000100000001000000010", 17963=>X"00000010000000100000001000000010", 17964=>X"00000010000000100000001000000010", 
17965=>X"00000010000000100000001000000010", 17966=>X"00000010000000100000001000000010", 17967=>X"00000010000000100000001000000010", 17968=>X"00000010000000100000001000000010", 17969=>X"00000010000000100000001000000010", 
17970=>X"00000010000000100000001000000010", 17971=>X"00000010000000100000001000000010", 17972=>X"00000010000000100000001000000010", 17973=>X"00000010000000100000001000000010", 17974=>X"00000010000000100000001000000010", 
17975=>X"00000010000000100000001000000010", 17976=>X"00000010000000100000001000000010", 17977=>X"00000010000000100000001000000010", 17978=>X"00000010000000100000001000000010", 17979=>X"00000010000000100000001000000010", 
17980=>X"00000010000000100000001000000010", 17981=>X"00000010000000100000001000000010", 17982=>X"00000010000000100000001000000010", 17983=>X"00000010000000100000001000000010", 17984=>X"00000010000000100000001000000010", 
17985=>X"00000010000000100000001000000010", 17986=>X"00000010000000100000001000000010", 17987=>X"00000010000000100000001000000010", 17988=>X"00000010000000100000001000000010", 17989=>X"00000010000000100000001000000010", 
17990=>X"00000010000000100000001000000010", 17991=>X"00000010000000100000001000000010", 17992=>X"00000010000000100000001000000010", 17993=>X"00000010000000100000001000000010", 17994=>X"00000010000000100000001000000010", 
17995=>X"00000010000000100000001000000010", 17996=>X"00000010000000100000001000000010", 17997=>X"00000010000000100000001000000010", 17998=>X"00000010000000100000001000000010", 17999=>X"00000010000000100000001000000010", 
18000=>X"00000010000000100000001000000010", 18001=>X"00000010000000100000001000000010", 18002=>X"00000010000000100000001000000010", 18003=>X"00000010000000100000001000000010", 18004=>X"00000010000000100000001000000010", 
18005=>X"00000010000000100000001000000010", 18006=>X"00000010000000100000001000000010", 18007=>X"00000010000000100000001000000010", 18008=>X"00000010000000100000001000000010", 18009=>X"00000010000000100000001000000010", 
18010=>X"00000010000000100000001000000010", 18011=>X"00000010000000100000001000000010", 18012=>X"00000010000000100000001000000010", 18013=>X"00000010000000100000001000000010", 18014=>X"00000010000000100000001000000010", 
18015=>X"00000010000000100000001000000010", 18016=>X"00000010000000100000001000000010", 18017=>X"00000010000000100000001000000010", 18018=>X"00000010000000100000001000000010", 18019=>X"00000010000000100000001000000010", 
18020=>X"00000010000000100000001000000010", 18021=>X"00000010000000100000001000000010", 18022=>X"00000010000000100000001000000010", 18023=>X"00000010000000100000001000000010", 18024=>X"00000010000000100000001000000010", 
18025=>X"00000010000000100000001000000010", 18026=>X"00000010000000100000001000000010", 18027=>X"00000010000000100000001000000010", 18028=>X"00000010000000100000001000000010", 18029=>X"00000010000000100000001000000010", 
18030=>X"00000010000000100000001000000010", 18031=>X"00000010000000100000001000000010", 18032=>X"00000010000000100000001000000010", 18033=>X"00000010000000100000001000000010", 18034=>X"00000010000000100000001000000010", 
18035=>X"00000010000000100000001000000010", 18036=>X"00000010000000100000001000000010", 18037=>X"00000010000000100000001000000010", 18038=>X"00000010000000100000001000000010", 18039=>X"00000010000000100000001000000010", 
18040=>X"00000010000000100000001000000010", 18041=>X"00000010000000100000001000000010", 18042=>X"00000010000000100000001000000010", 18043=>X"00000010000000100000001000000010", 18044=>X"00000010000000100000001000000010", 
18045=>X"00000010000000100000001000000010", 18046=>X"00000010000000100000001000000010", 18047=>X"00000010000000100000001000000010", 18048=>X"00000010000000100000001000000010", 18049=>X"00000010000000100000001000000010", 
18050=>X"00000010000000100000001000000010", 18051=>X"00000010000000100000001000000010", 18052=>X"00000010000000100000001000000010", 18053=>X"00000010000000100000001000000010", 18054=>X"00000010000000100000001000000010", 
18055=>X"00000010000000100000001000000010", 18056=>X"00000010000000100000001000000010", 18057=>X"00000010000000100000001000000010", 18058=>X"00000010000000100000001000000010", 18059=>X"00000010000000100000001000000010", 
18060=>X"00000010000000100000001000000010", 18061=>X"00000010000000100000001000000010", 18062=>X"00000010000000100000001000000010", 18063=>X"00000010000000100000001000000010", 18064=>X"00000010000000100000001000000010", 
18065=>X"00000010000000100000001000000010", 18066=>X"00000010000000100000001000000010", 18067=>X"00000010000000100000001000000010", 18068=>X"00000010000000100000001000000010", 18069=>X"00000010000000100000001000000010", 
18070=>X"00000010000000100000001000000010", 18071=>X"00000010000000100000001000000010", 18072=>X"00000010000000100000001000000010", 18073=>X"00000010000000100000001000000010", 18074=>X"00000010000000100000001000000010", 
18075=>X"00000010000000100000001000000010", 18076=>X"00000010000000100000001000000010", 18077=>X"00000010000000100000001000000010", 18078=>X"00000010000000100000001000000010", 18079=>X"00000010000000100000001000000010", 
18080=>X"00000010000000100000001000000010", 18081=>X"00000010000000100000001000000010", 18082=>X"00000010000000100000001000000010", 18083=>X"00000010000000100000001000000010", 18084=>X"00000010000000100000001000000010", 
18085=>X"00000010000000100000001000000010", 18086=>X"00000010000000100000001000000010", 18087=>X"00000010000000100000001000000010", 18088=>X"00000010000000100000001000000010", 18089=>X"00000010000000100000001000000010", 
18090=>X"00000010000000100000001000000010", 18091=>X"00000010000000100000001000000010", 18092=>X"00000010000000100000001000000010", 18093=>X"00000010000000100000001000000010", 18094=>X"00000010000000100000001000000010", 
18095=>X"00000010000000100000001000000010", 18096=>X"00000010000000100000001000000010", 18097=>X"00000010000000100000001000000010", 18098=>X"00000010000000100000001000000010", 18099=>X"00000010000000100000001000000010", 
18100=>X"00000010000000100000001000000010", 18101=>X"00000010000000100000001000000010", 18102=>X"00000010000000100000001000000010", 18103=>X"00000010000000100000001000000010", 18104=>X"00000010000000100000001000000010", 
18105=>X"00000010000000100000001000000010", 18106=>X"00000010000000100000001000000010", 18107=>X"00000010000000100000001000000010", 18108=>X"00000010000000100000001000000010", 18109=>X"00000010000000100000001000000010", 
18110=>X"00000010000000100000001000000010", 18111=>X"00000010000000100000001000000010", 18112=>X"00000010000000100000001000000010", 18113=>X"00000010000000100000001000000010", 18114=>X"00000010000000100000001000000010", 
18115=>X"00000010000000100000001000000010", 18116=>X"00000010000000100000001000000010", 18117=>X"00000010000000100000001000000010", 18118=>X"00000010000000100000001000000010", 18119=>X"00000010000000100000001000000010", 
18120=>X"00000010000000100000001000000010", 18121=>X"00000010000000100000001000000010", 18122=>X"00000010000000100000001000000010", 18123=>X"00000010000000100000001000000010", 18124=>X"00000010000000100000001000000010", 
18125=>X"00000010000000100000001000000010", 18126=>X"00000010000000100000001000000010", 18127=>X"00000010000000100000001000000010", 18128=>X"00000010000000100000001000000010", 18129=>X"00000010000000100000001000000010", 
18130=>X"00000010000000100000001000000010", 18131=>X"00000010000000100000001000000010", 18132=>X"00000010000000100000001000000010", 18133=>X"00000010000000100000001000000010", 18134=>X"00000010000000100000001000000010", 
18135=>X"00000010000000100000001000000010", 18136=>X"00000010000000100000001000000010", 18137=>X"00000010000000100000001000000010", 18138=>X"00000010000000100000001000000010", 18139=>X"00000010000000100000001000000010", 
18140=>X"00000010000000100000001000000010", 18141=>X"00000010000000100000001000000010", 18142=>X"00000010000000100000001000000010", 18143=>X"00000010000000100000001000000010", 18144=>X"00000010000000100000001000000010", 
18145=>X"00000010000000100000001000000010", 18146=>X"00000010000000100000001000000010", 18147=>X"00000010000000100000001000000010", 18148=>X"00000010000000100000001000000010", 18149=>X"00000010000000100000001000000010", 
18150=>X"00000010000000100000001000000010", 18151=>X"00000010000000100000001000000010", 18152=>X"00000010000000100000001000000010", 18153=>X"00000010000000100000001000000010", 18154=>X"00000010000000100000001000000010", 
18155=>X"00000010000000100000001000000010", 18156=>X"00000010000000100000001000000010", 18157=>X"00000010000000100000001000000010", 18158=>X"00000010000000100000001000000010", 18159=>X"00000010000000100000001000000010", 
18160=>X"00000010000000100000001000000010", 18161=>X"00000010000000100000001000000010", 18162=>X"00000010000000100000001000000010", 18163=>X"00000010000000100000001000000010", 18164=>X"00000010000000100000001000000010", 
18165=>X"00000010000000100000001000000010", 18166=>X"00000010000000100000001000000010", 18167=>X"00000010000000100000001000000010", 18168=>X"00000010000000100000001000000010", 18169=>X"00000010000000100000001000000010", 
18170=>X"00000010000000100000001000000010", 18171=>X"00000010000000100000001000000010", 18172=>X"00000010000000100000001000000010", 18173=>X"00000010000000100000001000000010", 18174=>X"00000010000000100000001000000010", 
18175=>X"00000010000000100000001000000010", 18176=>X"00000010000000100000001000000010", 18177=>X"00000010000000100000001000000010", 18178=>X"00000010000000100000001000000010", 18179=>X"00000010000000100000001000000010", 
18180=>X"00000010000000100000001000000010", 18181=>X"00000010000000100000001000000010", 18182=>X"00000010000000100000001000000010", 18183=>X"00000010000000100000001000000010", 18184=>X"00000010000000100000001000000010", 
18185=>X"00000010000000100000001000000010", 18186=>X"00000010000000100000001000000010", 18187=>X"00000010000000100000001000000010", 18188=>X"00000010000000100000001000000010", 18189=>X"00000010000000100000001000000010", 
18190=>X"00000010000000100000001000000010", 18191=>X"00000010000000100000001000000010", 18192=>X"00000010000000100000001000000010", 18193=>X"00000010000000100000001000000010", 18194=>X"00000010000000100000001000000010", 
18195=>X"00000010000000100000001000000010", 18196=>X"00000010000000100000001000000010", 18197=>X"00000010000000100000001000000010", 18198=>X"00000010000000100000001000000010", 18199=>X"00000010000000100000001000000010", 
18200=>X"00000010000000100000001000000010", 18201=>X"00000010000000100000001000000010", 18202=>X"00000010000000100000001000000010", 18203=>X"00000010000000100000001000000010", 18204=>X"00000010000000100000001000000010", 
18205=>X"00000010000000100000001000000010", 18206=>X"00000010000000100000001000000010", 18207=>X"00000010000000100000001000000010", 18208=>X"00000010000000100000001000000010", 18209=>X"00000010000000100000001000000010", 
18210=>X"00000010000000100000001000000010", 18211=>X"00000010000000100000001000000010", 18212=>X"00000010000000100000001000000010", 18213=>X"00000010000000100000001000000010", 18214=>X"00000010000000100000001000000010", 
18215=>X"00000010000000100000001000000010", 18216=>X"00000010000000100000001000000010", 18217=>X"00000010000000100000001000000010", 18218=>X"00000010000000100000001000000010", 18219=>X"00000010000000100000001000000010", 
18220=>X"00000010000000100000001000000010", 18221=>X"00000010000000100000001000000010", 18222=>X"00000010000000100000001000000010", 18223=>X"00000010000000100000001000000010", 18224=>X"00000010000000100000001000000010", 
18225=>X"00000010000000100000001000000010", 18226=>X"00000010000000100000001000000010", 18227=>X"00000010000000100000001000000010", 18228=>X"00000010000000100000001000000010", 18229=>X"00000010000000100000001000000010", 
18230=>X"00000010000000100000001000000010", 18231=>X"00000010000000100000001000000010", 18232=>X"00000010000000100000001000000010", 18233=>X"00000010000000100000001000000010", 18234=>X"00000010000000100000001000000010", 
18235=>X"00000010000000100000001000000010", 18236=>X"00000010000000100000001000000010", 18237=>X"00000010000000100000001000000010", 18238=>X"00000010000000100000001000000010", 18239=>X"00000010000000100000001000000010", 
18240=>X"00000010000000100000001000000010", 18241=>X"00000010000000100000001000000010", 18242=>X"00000010000000100000001000000010", 18243=>X"00000010000000100000001000000010", 18244=>X"00000010000000100000001000000010", 
18245=>X"00000010000000100000001000000010", 18246=>X"00000010000000100000001000000010", 18247=>X"00000010000000100000001000000010", 18248=>X"00000010000000100000001000000010", 18249=>X"00000010000000100000001000000010", 
18250=>X"00000010000000100000001000000010", 18251=>X"00000010000000100000001000000010", 18252=>X"00000010000000100000001000000010", 18253=>X"00000010000000100000001000000010", 18254=>X"00000010000000100000001000000010", 

-- OneDividedByDivision Constants
18255=>X"f4ffeefff4fff1fff4fff5fff4fff9ff",-- 8Sound samples
18256=>X"2b00300039003e004100490049005000"
);

begin

process(rst_n,clk,rd,wr,addr)
	variable regVal	:	std_logic_vector(127 downto 0);
	variable romWr : std_logic_vector (15 downto 0);	
begin
    
	data_out <= regVal;
	
    if rst_n='0' then
		regVal :=(others=>'0');
		ack <='0';
		
    elsif rising_edge(clk) then
		ack <='0';
		if cen='0' and (wr='0' or rd='0') then
            ack <='1'; --
            if unsigned(addr) <= MAX_ROWS then
                if wr='0' then
                    romWr := data_in;
                elsif rd='0' then
                    regVal := romRd(to_integer(unsigned(addr)));
                end if;
            end if;
            
       end if;--cen='0'		
	end if;
end process;
  
end Behavioral;
